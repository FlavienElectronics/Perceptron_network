-- VHDL Memory Module for Layer Weights: test_weights
-- Number of Neurons: 10
-- Number of Inputs per Neuron: 784
-- Data Width: 32 bits
-- Address Width: 10 bits
-- Expected Data Encoding: fixed_point
-- Res for 0x02000000 : 0x[]
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity test_weights is
    port(
        clk   : in  std_logic;
        addr  : in  std_logic_vector(9 downto 0); -- Same addr for all neurons within a layer
        dout  : out std_logic_vector(32*10-1 downto 0) -- DATA_WIDTH * N_NEURONS -> 320 bits
    );
end test_weights;

architecture rtl of test_weights is
    constant DATA_WIDTH : integer := 32;
    constant N_INPUTS  : integer := 784;
   type weight_array is array (0 to N_INPUTS-1) of std_logic_vector(DATA_WIDTH-1 downto 0);
    constant weights_n0 : weight_array := (
     x"FFCF3957", x"FF3ACB12", x"011DD0E0", x"FFC550EE", x"007434D5", x"FEFAC26C", x"00A86C6E", x"FFA512D5", x"FF217306", x"002AC7D9", x"008DBD5C", x"00FD30C3", x"FF4D45D4", x"FF6F848A", x"0037C086", x"004F57AE", x"00707C50", x"00A095D0", x"FFBDA889", x"00A28B37", x"00D7B5E1", x"FFB392F5", x"00D026EE", x"008EF1C5", x"0102103E", x"FF59BD42", x"FF6F868D", x"FFAB67FE", x"000ED750", x"00AF99E1", x"FF58FB5D", x"00927A20", x"FF97243E", x"00B0B9FE", x"FFF1E7DE", x"FEFEFF82", x"FF5DC1BD", x"FF2A28FA", x"008EE4CF", x"FF3B9324", x"FFE90F38", x"003D6CEE", x"FF5ADF56", x"0052D06D", x"FEE40E02", x"FF2E8965", x"FEF4F976", x"FFA5D843", x"FF93DC1E", x"0029429B", x"FFC9BACE", x"008985B4", x"010C3A68", x"0068F8D7", x"FF8CBC82", x"FEEE0A52", x"0069F84E", x"FF6F0B0D", x"0094E1B9", x"00C41585", x"0070D56F", x"01125680", x"01141CE0", x"003B811A", x"FF23A9E3", x"00F433D9", x"FF5BDF54", x"FF5699F9", x"00CAF9DC", x"00AA3BBE", x"000C8050", x"FFBD6249", x"FEB51266", x"FF8DFA49", x"00CAC040", x"00098E01", x"FFEE4ED1", x"FFABEB38", x"FF8D77C5", x"00A9690E", x"00109FC2", x"00BE0A32", x"FFCC371C", x"007FD3C0", x"0078C3C2", x"002EA797", x"00B7D756", x"00B87C7A", x"010E995A", x"00DAA9F4", x"FFA84A64", x"FEF03C5C", x"00102B73", x"FFB3A9F6", x"FF4F5EBA", x"FF6416C6", x"FF83671C", x"002DB3DB", x"FF8C2F7F", x"FEB31844", x"FE8EAB9C", x"FEA1A9CE", x"FE6B62AE", x"00069DBC", x"FFD8389D", x"00803C77", x"FFAF3D32", x"0016C22E", x"00589B7B", x"FEE90EF2", x"0019DAC1", x"FFEC6E0E", x"FF5BF7F9", x"FF1CFAB0", x"0102F954", x"00EE907B", x"0083D2B3", x"00FFBF02", x"FF56A668", x"FF7CD05E", x"FFF099E4", x"FF1F114D", x"FEF179A6", x"FE47E1E2", x"FFBDC706", x"FF3F2628", x"00418587", x"019673EC", x"FFCB0E25", x"FF8ED6A5", x"00502D7C", x"FF0ABA63", x"FF4493C1", x"0065863A", x"FF026BA3", x"FED7C24A", x"FF2BF033", x"FFA1AAC9", x"FF729BBB", x"FF681FFE", x"00762EC0", x"0031B80B", x"FFA22ECC", x"FF1C81A0", x"FF93D045", x"FF49BA86", x"FF322899", x"FE3F754C", x"FF32A41E", x"FDF878F0", x"FE221EF2", x"FE970246", x"00A275A5", x"009DBAB5", x"01988E0C", x"035D9988", x"03198088", x"02DE3AAC", x"0080DF37", x"000635C4", x"FFAEABC6", x"009A9B3E", x"FF80B56A", x"FE6DFCE2", x"FF85D32D", x"FEEE757A", x"FFB4E65B", x"FFAEB37B", x"00FD4493", x"005A9E00", x"FFCC185F", x"002A2170", x"FF876332", x"001E79BA", x"FFCBD67B", x"FF426FE0", x"FE350F2E", x"FFA3946D", x"FF127808", x"FF8717CB", x"015A6748", x"027E0CD0", x"03464844", x"03099DBC", x"02EF7C5C", x"044A86B8", x"0431E240", x"01160E0A", x"011AF556", x"FFEDFDF3", x"002F7EF5", x"FFBBEAEC", x"FEE2F2DE", x"FF73BB8A", x"0063DA0A", x"FFCC291D", x"FF0A4DEE", x"00E9D38C", x"FF691F35", x"FFD1860A", x"FFDAF04D", x"FF6D2AEC", x"FE0C2BF0", x"FF538060", x"FE24D77E", x"FE842746", x"FFEE52C7", x"FFA89695", x"0056A738", x"00FBE8BA", x"017476B8", x"02089EC4", x"03104790", x"0489ACA0", x"034CEDA0", x"0252C940", x"01AD8FA6", x"013B6298", x"01467F9A", x"FEF53F84", x"FF5EFA1A", x"FFF2B264", x"0073AF1B", x"FEF00B44", x"FF91A729", x"FF03C09C", x"FF3CF6DC", x"007EF2D4", x"FF698013", x"FFC493F0", x"FE5D5ED2", x"FF0DE878", x"FE5A9968", x"FFE9ADA0", x"FF58C5BF", x"00203677", x"0008A8E0", x"0162A602", x"02D6D3C0", x"02B9E4EC", x"026E8458", x"03B22818", x"03ED5738", x"024FFFF4", x"02F772DC", x"0161B1E0", x"01A24138", x"003E6F18", x"FECEFED0", x"FF6EEC88", x"003FB3CB", x"003F2527", x"FF72C225", x"011A9FA8", x"FFC5F3AA", x"FF19834E", x"FEF3E738", x"005B795C", x"FF31E988", x"FF213000", x"FEDE4BFC", x"FF5DA376", x"FF303662", x"FFC9F5E0", x"02204334", x"02B2AE28", x"0277AB10", x"0020ACC4", x"01D896C6", x"0148E324", x"03CFCB60", x"042290F8", x"0356D18C", x"02E9F288", x"03279488", x"01E378FA", x"009905F4", x"FEFFB812", x"005C5C88", x"FFA007C7", x"FFFAA673", x"FEFEC96E", x"FFA5300E", x"FF290D72", x"FF142240", x"FE9F62C6", x"FE913D96", x"FFE8DB32", x"007F286E", x"0105A0C6", x"010A6732", x"00D7F568", x"0093C33D", x"0177CC2C", x"007B6ADB", x"FDA08500", x"FEAE9928", x"00933A4C", x"01C73F2E", x"022832D4", x"04193330", x"03B99054", x"04AE6F78", x"02727CE0", x"017F0EC8", x"FEDBB92C", x"0104B2A6", x"FF832258", x"00AFFE32", x"0038C6EA", x"003BE520", x"FF95927D", x"FFE03807", x"FF1945B3", x"FF3DB04F", x"00315D76", x"0125D776", x"FFF261BF", x"016F7DE4", x"0166E378", x"01D0F0BA", x"FFF95E5D", x"FD72A188", x"FADAB8F0", x"FA283030", x"FCB5CB48", x"FEA6BB1A", x"02B965B8", x"021CACA8", x"04A9E008", x"0619BF78", x"04BE7B38", x"01D9EAAC", x"FEC3819C", x"010C5D36", x"FFCDA208", x"FEEE8AF0", x"011FAF40", x"FF7C53EA", x"FFB1B1D5", x"007EC8DC", x"FF4D8462", x"00592060", x"017FBA04", x"009122A0", x"016C7C4A", x"013A61CA", x"01C8056E", x"FF63D65C", x"FC5BA15C", x"F91374D8", x"F9392F38", x"F89CF948", x"F9386668", x"FE321022", x"00A71CC3", x"02A91E84", x"03970F4C", x"05AE05D0", x"05C1EF38", x"02B1BBF0", x"FF1E0DB7", x"0105C004", x"00167F5B", x"008CB750", x"00E39A78", x"00F2A6E5", x"FEEA6638", x"009A6126", x"000AA447", x"0211A434", x"0168B39E", x"0190397A", x"0259B650", x"02A08C04", x"00BE9101", x"FDEF8D98", x"FB62A6A0", x"F8BF8110", x"F7ACF420", x"F78CA170", x"F9E47A20", x"FC349A60", x"FF694B7C", x"01D72226", x"03068C08", x"0470C770", x"04C7DF88", x"01A03A74", x"000DB3F5", x"FFBA382F", x"002CE58F", x"00BE4C4B", x"FF9E9C6B", x"00E58711", x"00B59BC8", x"FEDB1528", x"00BA82F6", x"02033D9C", x"02A54958", x"0297828C", x"034B2F98", x"0262D1FC", x"FF07D8B7", x"FB694EC0", x"F81FB2F8", x"F7FD5830", x"F5F16590", x"F60B8760", x"F9F2E970", x"FC954F80", x"00443225", x"02309350", x"047A40B0", x"03BEF2E4", x"04EA7990", x"0304553C", x"FF8419D2", x"010A129C", x"00DB3E1F", x"00032E15", x"008CCD33", x"FF966F4F", x"FEC6FFF4", x"0038DC9B", x"02A0B8D0", x"02C7BD58", x"0488CD90", x"031E3084", x"05151B88", x"03627FDC", x"FE8188F8", x"F99ED418", x"F80F2640", x"F6804D40", x"F6A813E0", x"F81C9E00", x"FB9906B0", x"FD83D7BC", x"FFFF7AA7", x"01F079A8", x"02D259A8", x"048EA2F0", x"02E27114", x"01AE4C40", x"003EEB2E", x"FFADE64D", x"00C6DCA7", x"001FF70A", x"FEF169E2", x"FFDAC149", x"FF328653", x"002848C7", x"02778168", x"02D8184C", x"042CE798", x"048FD2A8", x"03CAE598", x"02D73478", x"FD503928", x"FA7AFEF8", x"F7D8E640", x"F5E708F0", x"F7B8CCF0", x"FA7AA0B8", x"FC19AA10", x"FEDDB6FE", x"022DA33C", x"0289F73C", x"019B2754", x"037EF2B0", x"026655B8", x"0000FE33", x"000BE2CF", x"0056557A", x"FFA75C95", x"0065C7E0", x"FF05B224", x"00C291FA", x"009C9546", x"00AE6279", x"02B03AA0", x"0453D9B0", x"03A62ED8", x"0475E130", x"041CB6C0", x"01358BA4", x"FCE6B4A4", x"FB4FACD0", x"F965D270", x"F729D9E0", x"F9ED8E48", x"FCB0CF4C", x"0016B394", x"01428F32", x"024F946C", x"00FB1B05", x"02720F38", x"0315ACBC", x"0078C4B8", x"FFA92AEA", x"002A3325", x"009A4006", x"FF70B7BE", x"00203372", x"FFFF6ED3", x"00405825", x"FEE166C6", x"00853FCD", x"02C8C570", x"029B530C", x"04460C10", x"04AB3BB0", x"0499CEC0", x"035089B8", x"FF2D18FF", x"FBC096A8", x"FB8E4320", x"FA3E6D08", x"FC1B91D0", x"FEB02950", x"FF7EAE07", x"0110CE8C", x"003D1770", x"00EC2183", x"013A6920", x"0169C118", x"FFC07251", x"FF07D3EA", x"007464DF", x"00F6DA5F", x"FEFB54AA", x"006C5DE0", x"FF2975A6", x"00043303", x"008C6A73", x"00A6CF5C", x"00A0BA7A", x"03643138", x"04183ED8", x"0427DC60", x"057BC980", x"02A72DC4", x"006DFD3A", x"FE122552", x"FD9D7FD4", x"FE10B416", x"FF08D201", x"FFB00014", x"007729FC", x"012116BC", x"FF637885", x"0026C33B", x"00A0622E", x"000F4029", x"00775757", x"FFEEB8C4", x"00B70592", x"FFE2B052", x"FF470134", x"00CEB785", x"002B954B", x"FFA0D3F4", x"FECD22B4", x"00112B5D", x"FFE6F4E0", x"0225E62C", x"02FEF18C", x"0260095C", x"0391FC8C", x"0339C858", x"03707208", x"01BB1A92", x"FFE1F432", x"00F2B16C", x"00589B72", x"FFEA13F8", x"0110E580", x"00659ECC", x"00D87348", x"FFF22A33", x"01067FDA", x"008C3510", x"007FB7C7", x"FEA9AF3E", x"00E00B72", x"FF041392", x"010649B6", x"FFF3E018", x"FEFC942A", x"00468A94", x"FF769E5E", x"FEC0B004", x"0024E1DC", x"01596F1E", x"02A32B14", x"021EC5B0", x"04632FB0", x"046F4320", x"03D90748", x"02B9F154", x"00EE35FB", x"00B1D1F5", x"013346D0", x"000120A0", x"FF8A9742", x"FF95052A", x"FEA4D33C", x"FF12F7C7", x"FF49C0B9", x"FF5A26C2", x"FF06539A", x"FFEC8806", x"FFCF56D8", x"00552A41", x"000D3A85", x"FF6DE5FD", x"FF9B43EF", x"FFF73AB0", x"FF1FAFDD", x"FFBC2D93", x"001245FC", x"0154DB8E", x"01AF802E", x"030C0680", x"032D9C5C", x"034A6618", x"0527A5C8", x"03A52F78", x"03E05C64", x"02BF88E4", x"01A5B59C", x"006398E6", x"00C2588F", x"FFB75375", x"FF5EED11", x"001C17DA", x"FE2A6C56", x"FFB3C518", x"0085B6E6", x"00B1E04A", x"FF1421F4", x"006854CE", x"FF595A11", x"FFF49170", x"FFC2F2F5", x"FF0A592D", x"FEDA24E0", x"FF0A0701", x"0056F2B8", x"0097FBEB", x"FF8DBB5D", x"00A594FB", x"01EF2BA2", x"01D7D1F4", x"04368888", x"04C0F758", x"03509B98", x"0138FB10", x"0115A74A", x"000517E0", x"FFCE4D6D", x"FE0A7E48", x"FDB781F8", x"FF79376D", x"FF6CE3AB", x"FF4F5D34", x"FF661F5A", x"FF6218ED", x"00EC284A", x"FFCD4AA3", x"00D3012C", x"010529EE", x"00250FD2", x"003D9D16", x"FFE92D17", x"00B94DEA", x"FED0E4C8", x"0031DA06", x"FF566195", x"FFF3047A", x"FF4D6376", x"FEE64376", x"FF3996DA", x"002BB963", x"FEC2C674", x"FE8D1C58", x"FEAA3F48", x"FE3267B6", x"FF08571B", x"FF8D4D06", x"FEF8B98C", x"00705201", x"FF1E8F9D", x"FF297191", x"FF6A05CE", x"FF3304D9", x"FF33A1E8", x"FEFB4EB2", x"FEFCB334", x"004C5C59", x"00B26D05", x"0112A4CA", x"00F8CC44", x"FFEAF9CB", x"0025B1EA", x"FF217AF2", x"001183C7", x"FE457D7E", x"FF9F0856", x"FEFC6DEE", x"FF086A95", x"FF07569E", x"FE29B514", x"FFB7CC6F", x"FF5CC0D0", x"FFA2E77C", x"FF2EBCDF", x"0003E0B6", x"0054057A", x"00369DCE", x"00ADCCB3", x"FFB36172", x"00B72456", x"0040F051", x"00B00615", x"011CF638", x"00423FC0", x"FF93683B", x"FFE2E3E9", x"00525E00", x"00314D52", x"FFAF4275", x"00DE1B00", x"009DF52A", x"FF2B7B82", x"FFB2D418", x"FF926BD5", x"FEE4C134", x"FFBDC800", x"FF3D0C18", x"FEFA02DC", x"FF2E1F51", x"FF2961D8", x"00B20531", x"00173287", x"00DC51C3", x"0029806C", x"0027557C", x"0065EBC4", x"00286AB8", x"FF185CE9", x"FF52EBDB", x"FFB9126F", x"000465F6", x"006E3745", x"0070A775", x"00E819D1", x"003B8F40", x"FF9C25B9", x"FF23F3E0", x"FF28EC23", x"FF4F713A", x"0055FC49", x"009A98F4", x"00FA31D2", x"FF9D9B0F", x"FFE20782", x"FF9B4A39", x"FFEBAA7C", x"004218D5", x"FFE1FD0A", x"FFF82A7F", x"0010CB5E", x"005D747F", x"FF9F467E", x"FF4CA807", x"004171EF", x"FFD66AA3", x"FF7A16E4", x"007ADE82", x"0002A742", x"FFD570F3", x"FF725EF4"
--  -0.005954, -0.024073, 0.034890, -0.007164, 0.014185, -0.031890, 0.020560, -0.011099, -0.027167, 0.005222, 0.017302, 0.030907, -0.021817, -0.017637, 0.006806, 0.009685, 0.013731, 0.019603, -0.008098, 0.019842, 0.026332, -0.009329, 0.025409, 0.017449, 0.031502, -0.020295, -0.017636, -0.010326, 0.001812, 0.021436, -0.020388, 0.017880, -0.012800, 0.021573, -0.001720, -0.031372, -0.019805, -0.026104, 0.017443, -0.023978, -0.002800, 0.007498, -0.020157, 0.010109, -0.034661, -0.025569, -0.032596, -0.011005, -0.013201, 0.005037, -0.006625, 0.016787, 0.032743, 0.012814, -0.014070, -0.033442, 0.012936, -0.017695, 0.018174, 0.023936, 0.013774, 0.033489, 0.033705, 0.007264, -0.026897, 0.029810, -0.020035, -0.020679, 0.024777, 0.020780, 0.001526, -0.008132, -0.040397, -0.013919, 0.024750, 0.001166, -0.002160, -0.010264, -0.013981, 0.020680, 0.002029, 0.023198, -0.006321, 0.015604, 0.014742, 0.005695, 0.022442, 0.022520, 0.033032, 0.026692, -0.010707, -0.033174, 0.001974, -0.009318, -0.021561, -0.019032, -0.015210, 0.005579, -0.014138, -0.040638, -0.045084, -0.042766, -0.049391, 0.000808, -0.004856, 0.015654, -0.009859, 0.002778, 0.010816, -0.034050, 0.003156, -0.002389, -0.020023, -0.027712, 0.031613, 0.029122, 0.016092, 0.031219, -0.020673, -0.016014, -0.001880, -0.027458, -0.033023, -0.053725, -0.008084, -0.023541, 0.007998, 0.049616, -0.006463, -0.013814, 0.009787, -0.029940, -0.022879, 0.012393, -0.030955, -0.036162, -0.025886, -0.011515, -0.017260, -0.018539, 0.014427, 0.006069, -0.011452, -0.027770, -0.013206, -0.022250, -0.025127, -0.054754, -0.025068, -0.063419, -0.058335, -0.044066, 0.019831, 0.019254, 0.049872, 0.105176, 0.096863, 0.089628, 0.015731, 0.000758, -0.009928, 0.018873, -0.015538, -0.049074, -0.014914, -0.033391, -0.009168, -0.009924, 0.030916, 0.011062, -0.006336, 0.005143, -0.014723, 0.003720, -0.006367, -0.023140, -0.056023, -0.011282, -0.028995, -0.014759, 0.042286, 0.077887, 0.102329, 0.094924, 0.091734, 0.134097, 0.131089, 0.033942, 0.034541, -0.002198, 0.005798, -0.008311, -0.034796, -0.017122, 0.012189, -0.006328, -0.029992, 0.028543, -0.018418, -0.005673, -0.004524, -0.017924, -0.061014, -0.021057, -0.058003, -0.046368, -0.002158, -0.010670, 0.010578, 0.030751, 0.045467, 0.063552, 0.095737, 0.141806, 0.103141, 0.072606, 0.052437, 0.038499, 0.039856, -0.032562, -0.019656, -0.001624, 0.014122, -0.033198, -0.013470, -0.030792, -0.023808, 0.015497, -0.018372, -0.007254, -0.051102, -0.029552, -0.051441, -0.002725, -0.020414, 0.003932, 0.001057, 0.043292, 0.088724, 0.085192, 0.075991, 0.115498, 0.122722, 0.072266, 0.092706, 0.043176, 0.051056, 0.007621, -0.037232, -0.017709, 0.007776, 0.007708, -0.017241, 0.034500, -0.007086, -0.028136, -0.032727, 0.011166, -0.025157, -0.027199, -0.035364, -0.019820, -0.025365, -0.006597, 0.066438, 0.084312, 0.077108, 0.003989, 0.057689, 0.040147, 0.119116, 0.129220, 0.104348, 0.091058, 0.098582, 0.059018, 0.018680, -0.031284, 0.011275, -0.011715, -0.000653, -0.031398, -0.011085, -0.026239, -0.028792, -0.043044, -0.044770, -0.002825, 0.015522, 0.031937, 0.032520, 0.026362, 0.018037, 0.045874, 0.015066, -0.074155, -0.041187, 0.017972, 0.055572, 0.067407, 0.128076, 0.116402, 0.146293, 0.076476, 0.046760, -0.035678, 0.031823, -0.015242, 0.021484, 0.006931, 0.007311, -0.012992, -0.003880, -0.028165, -0.023720, 0.006026, 0.035869, -0.001662, 0.044860, 0.043810, 0.056755, -0.000809, -0.079757, -0.160800, -0.182594, -0.102808, -0.042147, 0.085132, 0.066000, 0.145737, 0.190643, 0.148252, 0.057851, -0.038634, 0.032759, -0.006148, -0.033381, 0.035118, -0.016073, -0.009559, 0.015477, -0.021787, 0.010880, 0.046842, 0.017717, 0.044493, 0.038377, 0.055667, -0.019063, -0.113815, -0.216375, -0.211769, -0.230838, -0.211865, -0.056389, 0.020399, 0.083144, 0.112190, 0.177493, 0.179924, 0.084196, -0.027581, 0.031952, 0.002746, 0.017177, 0.027784, 0.029621, -0.033887, 0.018845, 0.001299, 0.064653, 0.044031, 0.048856, 0.073451, 0.082098, 0.023263, -0.064508, -0.144208, -0.226623, -0.260137, -0.264083, -0.190860, -0.118579, -0.018397, 0.057511, 0.094549, 0.138767, 0.149399, 0.050809, 0.001673, -0.008518, 0.005481, 0.023230, -0.011888, 0.028019, 0.022169, -0.035757, 0.022768, 0.062896, 0.082677, 0.080995, 0.102928, 0.074563, -0.030292, -0.143395, -0.246130, -0.250324, -0.314283, -0.311093, -0.189098, -0.106774, 0.008325, 0.068430, 0.139923, 0.117059, 0.153622, 0.094279, -0.015124, 0.032480, 0.026763, 0.000388, 0.017188, -0.012886, -0.038208, 0.006941, 0.082119, 0.086882, 0.141700, 0.097435, 0.158827, 0.105774, -0.046688, -0.199362, -0.248151, -0.296838, -0.291983, -0.246507, -0.137570, -0.077656, -0.000064, 0.060605, 0.088178, 0.142412, 0.090142, 0.052527, 0.007681, -0.010022, 0.024275, 0.003902, -0.033031, -0.004547, -0.025082, 0.004918, 0.077088, 0.088879, 0.130482, 0.142557, 0.118518, 0.088770, -0.083957, -0.172486, -0.254773, -0.315547, -0.258691, -0.172531, -0.121867, -0.035435, 0.068071, 0.079342, 0.050190, 0.109247, 0.074992, 0.000121, 0.001451, 0.010539, -0.010820, 0.012424, -0.030555, 0.023751, 0.019114, 0.021287, 0.084012, 0.135236, 0.114036, 0.139390, 0.128505, 0.037786, -0.096838, -0.146524, -0.206321, -0.276141, -0.189751, -0.103417, 0.002771, 0.039375, 0.072214, 0.030653, 0.076423, 0.096396, 0.014742, -0.010600, 0.005151, 0.018829, -0.017491, 0.003931, -0.000069, 0.007855, -0.034985, 0.016266, 0.087008, 0.081460, 0.133551, 0.145902, 0.143775, 0.103581, -0.025745, -0.132741, -0.138884, -0.179880, -0.121635, -0.040996, -0.015786, 0.033302, 0.007457, 0.028825, 0.038380, 0.044159, -0.007758, -0.030294, 0.014208, 0.030133, -0.031820, 0.013228, -0.026189, 0.000513, 0.017141, 0.020363, 0.019620, 0.105981, 0.127960, 0.129866, 0.171361, 0.082908, 0.013426, -0.060285, -0.074524, -0.060461, -0.030173, -0.009766, 0.014546, 0.035289, -0.019108, 0.004732, 0.019578, 0.001862, 0.014568, -0.002109, 0.022342, -0.003578, -0.022582, 0.025234, 0.005320, -0.011618, -0.037459, 0.002096, -0.003057, 0.067126, 0.093621, 0.074223, 0.111571, 0.100804, 0.107476, 0.054090, -0.003668, 0.029626, 0.010816, -0.002676, 0.033313, 0.012405, 0.026422, -0.001689, 0.032043, 0.017115, 0.015591, -0.041787, 0.027349, -0.030752, 0.032018, -0.001480, -0.031668, 0.008611, -0.016770, -0.038979, 0.004502, 0.042167, 0.082418, 0.066256, 0.137108, 0.138582, 0.120243, 0.085198, 0.029078, 0.021707, 0.037509, 0.000138, -0.014332, -0.013059, -0.042380, -0.028935, -0.022247, -0.020245, -0.030478, -0.002377, -0.005940, 0.010396, 0.001615, -0.017835, -0.012297, -0.001071, -0.027382, -0.008279, 0.002231, 0.041609, 0.052673, 0.095218, 0.099318, 0.102832, 0.161090, 0.113914, 0.121138, 0.085881, 0.051478, 0.012158, 0.023724, -0.008871, -0.019662, 0.003429, -0.057321, -0.009305, 0.016323, 0.021713, -0.028792, 0.012736, -0.020343, -0.001395, -0.007453, -0.029987, -0.035871, -0.030026, 0.010614, 0.018553, -0.013949, 0.020213, 0.060446, 0.057595, 0.131657, 0.148555, 0.103590, 0.038206, 0.033893, 0.000622, -0.006067, -0.061219, -0.071349, -0.016453, -0.017958, -0.021562, -0.018784, -0.019275, 0.028828, -0.006190, 0.025757, 0.031880, 0.004524, 0.007521, -0.002786, 0.022620, -0.037000, 0.006085, -0.020705, -0.001585, -0.021803, -0.034392, -0.024220, 0.005337, -0.038724, -0.045275, -0.041718, -0.056347, -0.030232, -0.014001, -0.032138, 0.013711, -0.027519, -0.026191, -0.018308, -0.025022, -0.024947, -0.031823, -0.031653, 0.009321, 0.021781, 0.033526, 0.030371, -0.002566, 0.004601, -0.027163, 0.002138, -0.054017, -0.011837, -0.031686, -0.030223, -0.030354, -0.057409, -0.008814, -0.019928, -0.011364, -0.025545, 0.000473, 0.010257, 0.006667, 0.021216, -0.009353, 0.022356, 0.007927, 0.021487, 0.034785, 0.008087, -0.013256, -0.003553, 0.010055, 0.006018, -0.009856, 0.027112, 0.019282, -0.025942, -0.009420, -0.013376, -0.034576, -0.008083, -0.023798, -0.031981, -0.025620, -0.026198, 0.021731, 0.002832, 0.026894, 0.005066, 0.004802, 0.012442, 0.004934, -0.028276, -0.021128, -0.008658, 0.000537, 0.013454, 0.013752, 0.028333, 0.007270, -0.012189, -0.026861, -0.026255, -0.021552, 0.010496, 0.018872, 0.030541, -0.012011, -0.003659, -0.012294, -0.002482, 0.008068, -0.003664, -0.000956, 0.002050, 0.011408, -0.011807, -0.021893, 0.007989, -0.005076, -0.016347, 0.014999, 0.000324, -0.005195, -0.017289
--  Sum of weights (converted): 000000005AF884A0
    );

    constant weights_n1 : weight_array := (
     x"FFD981F0", x"FF07381B", x"00428EA2", x"000463F9", x"00B18B03", x"0012E436", x"00176449", x"004FB345", x"00DEA0EC", x"FF75BE3D", x"00AEAAAA", x"00478D3E", x"FF3CCA6B", x"00656D51", x"FF501DA5", x"FFA3E2FC", x"FF748A52", x"FF38F5A2", x"00E66BC1", x"FEFA7E58", x"00924A45", x"FEF8AEA6", x"FFDC646E", x"00117319", x"00CFFDFC", x"FF961ECB", x"005435C9", x"002D5230", x"00AC2505", x"001164D2", x"006D8D42", x"FF4F42A2", x"FF34AFCD", x"0104B290", x"FF2AC0C2", x"FFCDEB3D", x"FFDA833A", x"011BD0CE", x"FFBEFEF7", x"FF1F2E16", x"FFB3B2B9", x"00944590", x"0075B2A9", x"00F68FED", x"FFC00BD3", x"0086480F", x"FEEAE7C4", x"00703AFE", x"0085A5D5", x"00BC47D1", x"FF581A02", x"FFB1E113", x"0046C820", x"FF30182D", x"FF1743D6", x"FEE688A4", x"00105509", x"00B5AEEE", x"004B265C", x"0011CF8B", x"0065C3F8", x"FF481590", x"001E6484", x"FFB51769", x"FF679010", x"00EECB2C", x"FF0A0BAA", x"0015B8FB", x"FEEC5184", x"FFEFBD38", x"FF7E5F00", x"006F3DE8", x"FF54F31E", x"009DA854", x"FEEE295E", x"008FA8FA", x"FF098673", x"008B40B9", x"FF7AC346", x"FFFB69BE", x"FFC92BC1", x"00BDA1BC", x"005FE23B", x"FEFE2F4C", x"001AE630", x"FF362A7D", x"00DACCF0", x"00300349", x"FFB49E84", x"FF693766", x"00607910", x"FF4021ED", x"005F1491", x"00526BAD", x"003CA6E7", x"FFB49B7D", x"FE6677C6", x"0055D94A", x"FF379DFB", x"FF4AE3EC", x"FF58F0EC", x"00164A34", x"001B38DC", x"FF82C3E2", x"000EDADA", x"FEA714D0", x"FFDD9321", x"FEEA566E", x"0058259C", x"FF2D397C", x"FF96B872", x"00CC843E", x"01179BFC", x"FF50583B", x"FF5DE6C9", x"002427E4", x"007289EC", x"FFCBBF14", x"FF8CF66F", x"FEF94FA0", x"FFF802E6", x"004F8968", x"FE93824C", x"FFFA4D95", x"00DBA772", x"020E2CD4", x"011CB224", x"00EC9880", x"010F4C84", x"00A78034", x"01682E1A", x"00E3F228", x"020F3878", x"022849C4", x"FFF1F1A1", x"006F2AFD", x"FFAD1394", x"00AD0370", x"FF79CE57", x"0013C8C2", x"00AF0C73", x"FEF3F868", x"FF096DEB", x"FF6BDCE1", x"00BA08B8", x"00AF8969", x"FEEE98E2", x"FF8F0038", x"FE31524A", x"FDCDB0C0", x"FF4B4BBA", x"FF84BA97", x"0006CAED", x"01D46B66", x"01C6DF64", x"011146DC", x"FF4CDA12", x"FED8EB9E", x"01399220", x"02013300", x"0329DE98", x"01E68E8C", x"01C62604", x"012A20B4", x"009B567E", x"002566E6", x"0117D4DC", x"FFFE7637", x"003E49A0", x"0115F9FC", x"011B126A", x"FF85686A", x"00FA9AAF", x"002E23DF", x"FF4622BB", x"FFCB0003", x"FD635B54", x"FDE95BA0", x"FE166C6E", x"FCDCEA34", x"FE45F770", x"FEFF7230", x"FFC70EFC", x"FD912488", x"FD1DEFB0", x"FE22FE70", x"006C834E", x"01E4D464", x"02882550", x"01AADEB4", x"FF8A0E4B", x"FED04134", x"FF9C99E7", x"00C92161", x"0001B234", x"FFE385C0", x"FF396BB9", x"FF6E98B5", x"FF1D865D", x"00E338BD", x"FFB50463", x"FE8FAB14", x"FF1D50A5", x"FE602EA0", x"FD188478", x"FCB95688", x"FC69C364", x"FB0418A8", x"FCB4C658", x"FEFD2710", x"FE174EF6", x"FD087254", x"FE35726C", x"FDA3B914", x"FEA88448", x"FFFD020E", x"FF552ECF", x"005DF340", x"FEBCD4A4", x"FE2DDBD8", x"FE232A5E", x"002AC704", x"FFC053E1", x"FFDE0E04", x"FFB3BE5F", x"FF7287BC", x"0031C3B0", x"00D65169", x"FF2FB9BD", x"FF81EBD5", x"FDF17100", x"FD798C10", x"FDFAA614", x"FBF240D8", x"FC4ACBA4", x"FB349110", x"FC6171A8", x"FE8BBCDE", x"01970AEA", x"FFC61C6F", x"FFFFA063", x"FFA14B36", x"FFC3CE85", x"FFAADB39", x"FDFA2FF8", x"FE689728", x"FCCD0A3C", x"FDAAC6BC", x"FF7CB54A", x"FFB4A68F", x"FFC09718", x"FFBA4F11", x"FF4D29DA", x"00B1CBA1", x"FFF2FB2C", x"FFE93499", x"001BBDB7", x"00480D1D", x"FE4756C4", x"FDC56A44", x"FDEF5D44", x"FCD2DE40", x"FAE1A550", x"FA53A770", x"FD45123C", x"010062BE", x"03DB7BE4", x"05653A88", x"016B4E12", x"00B92C3C", x"FE313B46", x"FE4C9312", x"FDB66A8C", x"FD311078", x"FE4E670A", x"FD576DB4", x"FDC90028", x"FE66DB74", x"00A72679", x"0064C917", x"FF2983A9", x"008DFD74", x"0107A24C", x"FED2A140", x"00AEDFC2", x"FFB0E4A7", x"FF13CDDC", x"FF64CD6B", x"FE8C4BB0", x"FCF9AA14", x"FC98364C", x"FBD63C10", x"FD31AD64", x"00890037", x"07610120", x"07818E68", x"043AB960", x"00084810", x"FDE85DDC", x"FC0E6900", x"FBD5CB18", x"FE0863FE", x"FE96F43E", x"FF4E30D6", x"FEE910B4", x"FF8AB05B", x"FFA981FA", x"00C88CB5", x"FF81A038", x"00B815B9", x"00C79BD8", x"FEEB57B0", x"FFE84F08", x"FF6C226D", x"FE85F4AC", x"FF07C44F", x"FD846BC0", x"FD750258", x"FAA743A0", x"FB2221B8", x"FB4F1108", x"020B2B18", x"0A8A3B00", x"0B8D9BC0", x"0428EBC8", x"FDC9E6B0", x"FD492DA8", x"FBF4E1C0", x"FD3E60A4", x"FD32D5E8", x"FE83316A", x"001A8A55", x"FE99FB48", x"FECB2010", x"002E950A", x"00285020", x"FFCA7A64", x"00FF4F3C", x"FF4E3A1C", x"FF492A04", x"FF13EAE5", x"FF740BBA", x"FEFD6DDA", x"FF620D5F", x"FDA6C0B8", x"FCB400B0", x"FA3147E0", x"FA766550", x"FC666F4C", x"02E26678", x"0CC07750", x"099FB670", x"024E1100", x"FC5FFEFC", x"FBBBCF80", x"FDDB6EC4", x"FCC66020", x"FF8EF4D6", x"FF49BB21", x"0073AA1C", x"FF30E697", x"00B012B7", x"001EF254", x"001669D3", x"00C7C0F5", x"FEE9D568", x"FF137193", x"01180C80", x"FF41C2C0", x"FED9EA8C", x"FF35FC9F", x"FE38F466", x"FD7B6C60", x"FB3817D8", x"FA58C8D0", x"F7B7A2E0", x"FB3C0850", x"06A07A50", x"0DAC64B0", x"091B06A0", x"FFB0B30A", x"FB27D860", x"FB4550C0", x"FC6DB138", x"FD531734", x"FE34EC6E", x"005480F2", x"FF4A3344", x"001BC212", x"00B50870", x"FFE35847", x"FF61E198", x"FF39C500", x"FF9427EB", x"0068268C", x"FF09A981", x"FFCEF1CF", x"0014E200", x"0018B789", x"FED08616", x"FDB67F20", x"FC8D5E58", x"FA447AE0", x"F9278788", x"FC712EF4", x"07154330", x"0C3EA7A0", x"069DA518", x"FCDE27B4", x"F9B9A000", x"FB95B2B0", x"FD7BFB90", x"FD7095EC", x"FD924B34", x"FE7D8FC4", x"FEDAFC1E", x"0054EF2B", x"FF2950D7", x"FFE01CAA", x"FFC1E42C", x"FF4E6D7A", x"0084990E", x"FF870DBE", x"FFEED447", x"FF1D3F2E", x"FF6F4177", x"FF242C3B", x"FE4642FA", x"FCF1A1D8", x"FC2934A0", x"F9F2F9F8", x"FA385D88", x"FF1CA132", x"08E41D50", x"0A850970", x"04D57498", x"FA517850", x"F8E2D208", x"FB16B9C8", x"FCC2A424", x"FD8444C4", x"FF35B439", x"FE3EF242", x"FFB8FF51", x"FF9EE3DF", x"FEF0CF3C", x"FF86C3BA", x"0049B16D", x"0037E3B9", x"00D4BB2A", x"00C4F1D5", x"FF57F013", x"FF5C8E1F", x"FF238534", x"FDD140B8", x"FD9F4458", x"FC302E7C", x"FC845ADC", x"FCACE04C", x"FDBF5990", x"016B7FDE", x"08859EE0", x"0976AF90", x"01777FFE", x"FA62E7B8", x"F9B1A4B0", x"FBFB9E20", x"FCEF3DB4", x"FDC7F634", x"FE20FD96", x"FF64D5F8", x"FFA69F22", x"FE86E608", x"FF1D24F8", x"FFFEC2C4", x"006E40EE", x"008E563C", x"FF522E8A", x"FEDB8192", x"FFE366F8", x"FFA13BB0", x"FF6576FF", x"FDC91580", x"FE50B7C2", x"FD10B5F8", x"FDB70118", x"FD5B1954", x"0099DD22", x"043959A8", x"081A7D80", x"07A1BEF8", x"FEAE005C", x"FBD56900", x"FA2C8AA0", x"FB412780", x"FD180804", x"FDB379CC", x"FECA38A4", x"FF847A85", x"FE4031BC", x"00381B24", x"FF926AAF", x"FFAF80B7", x"0039FE32", x"00E4C6FE", x"FF60F047", x"FF3719BE", x"009FF650", x"FF187168", x"FF1A5E7C", x"FD5FE6A8", x"FD5786D4", x"FE1C2ECE", x"FD95AE94", x"FF3111FC", x"02512388", x"047C2DF8", x"062EED90", x"0367A180", x"00595643", x"FBBA2E50", x"FAD75CA8", x"FB4E0540", x"FCB13850", x"FE580A34", x"FE4BC392", x"FFB42045", x"FF0749C1", x"FF509B14", x"0076EFF3", x"FFF24B6D", x"FFC6620D", x"0061CF63", x"00E69E16", x"00430AE4", x"00ADF4CD", x"0049533D", x"FEE0E862", x"FDE8A24C", x"FD88606C", x"FDF3C630", x"003E4188", x"01A8D232", x"025A8964", x"0292ECB8", x"04708E88", x"0156C46E", x"005882C1", x"FDA658BC", x"FCE6FA54", x"FC9A1C78", x"FCA4AEB8", x"FEDB0564", x"FDFEFC1C", x"FF2EA264", x"FFF04418", x"FE9368E8", x"FFF789D9", x"FF949AE9", x"00D03447", x"FF45B826", x"00B16353", x"00AF2069", x"007D06DF", x"00AAA233", x"FF0A2259", x"FD4BEF00", x"FF1412BB", x"FF293842", x"0041C04E", x"FFE6ED29", x"00B19B79", x"FFC2C076", x"019A70CA", x"017B8E3C", x"006CCE28", x"FF13C79C", x"FCE51E8C", x"FD246D70", x"FD7A9FD8", x"FDD6FD48", x"FF96FF4E", x"FF732628", x"005B6FBC", x"FFA7F915", x"FEE76A8C", x"FFA89393", x"00CDB735", x"00B229EA", x"005A86E8", x"FFA3808E", x"FEDA1304", x"FF331208", x"0065BE5D", x"FF61598D", x"00824AB5", x"00D91E58", x"006C8A2A", x"01310FD8", x"FEA157B8", x"FDDF1A94", x"FDEC1244", x"FEB3674E", x"0078DA37", x"0000FEC4", x"FE5E835A", x"FF34C830", x"FD6D1A0C", x"FDA11F98", x"FE58F0BE", x"FED77408", x"FF6B4D9D", x"FF9884A0", x"007DB893", x"FEFD1270", x"002B1497", x"00051C20", x"004D495A", x"011E8DAA", x"00A73783", x"FF63ECF8", x"FFB8FEB3", x"00C916C4", x"00DE82CC", x"020E12E0", x"013F181A", x"008998D1", x"FDE130B4", x"FC2A7C18", x"FD85C45C", x"002BD592", x"012BEF82", x"020B08F4", x"FF7B97C7", x"000C48AE", x"FE61370E", x"FE365060", x"FF19EA80", x"0008F787", x"008AD94E", x"0031F0E7", x"FFE61DA2", x"FFF02E62", x"FF8965A2", x"FFE5BED3", x"FFEBC8FC", x"00F82B94", x"00A1081D", x"FF2B0B10", x"00B25A0E", x"00AEB4FC", x"019709AC", x"00DC0227", x"01586478", x"FE6E1F3C", x"FE927A30", x"FE069026", x"FD72CEF4", x"FF0D850C", x"01B29DA8", x"01499F30", x"011D722A", x"FEF6DCA6", x"0004BE69", x"FE9C5D82", x"FF0C4F0C", x"FF2BACB5", x"006AB79C", x"FFEE8FAF", x"FEE6F108", x"FF59FB73", x"FF789ACD", x"FEF08B26", x"0025767D", x"006831AD", x"FFC50A1D", x"FF84275E", x"0024D149", x"FF566FD0", x"FF47B488", x"FF72BCAB", x"FFD44C05", x"FD6B6FD0", x"FD9D6B3C", x"FC913F80", x"FD2CB984", x"FD2BAA10", x"FFE0D691", x"00539311", x"FF82C491", x"005C7F34", x"00B185EE", x"0061DEBF", x"007D394B", x"FED658DA", x"FEE2EE62", x"FF1C6ADA", x"005C7BCF", x"FF03229C", x"FF20AACB", x"FF723096", x"FEF25758", x"00006448", x"00298266", x"FF4DD446", x"00AB4598", x"FF613D38", x"FF3A6D06", x"0021500D", x"FFDFEB29", x"FE50CB02", x"FD855C58", x"FDD44704", x"FE8BD374", x"FF450C78", x"FF676FA5", x"FEC01E36", x"FE83923A", x"FECB723A", x"FF8379FF", x"FFF1F0B2", x"FF735B3F", x"FF139963", x"001C8D01", x"FF16F68A", x"FF1F518B", x"FF122619", x"FFB0B88E", x"01026A86", x"00725F30", x"FFDD4F63", x"003C198D", x"007274B0", x"FFFD0BFF", x"FF0883B3", x"FF33DE35", x"FF129848", x"FFC2C401", x"FEA916DA", x"FF736C4D", x"FF366A6C", x"00B1CA5B", x"009340EB", x"006DAE1F", x"FFE6B829", x"FF87923E", x"003C1028", x"FF2D5A6D", x"FF7E46A6", x"FFC27196", x"FFBA409E", x"FEEA8586", x"00744673", x"00F0E50A", x"FF5EA019", x"004EDE0E", x"FFDE11B9", x"FFF55447", x"00110DD2", x"00FD898C", x"00272DB5", x"FF46A5BA", x"FF962048", x"008E2EF1", x"005A2954", x"0003F410", x"FFD594C1", x"FF8B4349", x"FF93C9BF", x"FF6091FC", x"002ACEE5", x"004DDDC8", x"00DBBFAF", x"FFB9B7DA", x"0011E72D", x"00BC568E", x"007EB9F0", x"002568B9", x"0059A793", x"000F2BD9", x"FF0508DD", x"000B4769", x"FFC00CD0", x"0108051A"
--  -0.004699, -0.030369, 0.008125, 0.000536, 0.021673, 0.002306, 0.002855, 0.009729, 0.027176, -0.016877, 0.021322, 0.008734, -0.023829, 0.012381, -0.021470, -0.011244, -0.017024, -0.024297, 0.028128, -0.031922, 0.017858, -0.032143, -0.004347, 0.002130, 0.025390, -0.012925, 0.010280, 0.005532, 0.021014, 0.002123, 0.013373, -0.021575, -0.024819, 0.031823, -0.026031, -0.006113, -0.004576, 0.034645, -0.007935, -0.027444, -0.009314, 0.018100, 0.014367, 0.030098, -0.007807, 0.016392, -0.033825, 0.013700, 0.016314, 0.022983, -0.020495, -0.009536, 0.008640, -0.025379, -0.028410, -0.034359, 0.001994, 0.022178, 0.009174, 0.002174, 0.012423, -0.022451, 0.003710, -0.009144, -0.018608, 0.029150, -0.030024, 0.002652, -0.033653, -0.001985, -0.015824, 0.013579, -0.020880, 0.019245, -0.033428, 0.017537, -0.030087, 0.016999, -0.016264, -0.000560, -0.006693, 0.023148, 0.011705, -0.031472, 0.003284, -0.024638, 0.026709, 0.005861, -0.009202, -0.018406, 0.011776, -0.023421, 0.011606, 0.010061, 0.007404, -0.009203, -0.049992, 0.010480, -0.024461, -0.022108, -0.020393, 0.002721, 0.003323, -0.015287, 0.001813, -0.042104, -0.004202, -0.033894, 0.010760, -0.025729, -0.012852, 0.024965, 0.034132, -0.021442, -0.019787, 0.004414, 0.013982, -0.006379, -0.014043, -0.032067, -0.000975, 0.009709, -0.044494, -0.000695, 0.026813, 0.064230, 0.034753, 0.028881, 0.033118, 0.020447, 0.043967, 0.027825, 0.064358, 0.067418, -0.001716, 0.013570, -0.010123, 0.021120, -0.016381, 0.002415, 0.021368, -0.032718, -0.030099, -0.018083, 0.022709, 0.021428, -0.033374, -0.013794, -0.056479, -0.068641, -0.022059, -0.015048, 0.000829, 0.057180, 0.055526, 0.033359, -0.021869, -0.036020, 0.038278, 0.062646, 0.098861, 0.059394, 0.055438, 0.036393, 0.018962, 0.004566, 0.034159, -0.000188, 0.007603, 0.033933, 0.034555, -0.014965, 0.030591, 0.005632, -0.022689, -0.006470, -0.081621, -0.065264, -0.059763, -0.098033, -0.053959, -0.031318, -0.006951, -0.076032, -0.090096, -0.058228, 0.013246, 0.059183, 0.079119, 0.052108, -0.014397, -0.037078, -0.012134, 0.024552, 0.000207, -0.003476, -0.024241, -0.017749, -0.027646, 0.027737, -0.009153, -0.044962, -0.027672, -0.050759, -0.090757, -0.102376, -0.112089, -0.155750, -0.102933, -0.031598, -0.059655, -0.092719, -0.055976, -0.073764, -0.041929, -0.000365, -0.020852, 0.011469, -0.039449, -0.056902, -0.058207, 0.005222, -0.007773, -0.004144, -0.009309, -0.017269, 0.006075, 0.026162, -0.025424, -0.015390, -0.064277, -0.078913, -0.063153, -0.126678, -0.115870, -0.149833, -0.113105, -0.045442, 0.049688, -0.007067, -0.000046, -0.011561, -0.007348, -0.010394, -0.063210, -0.049733, -0.099971, -0.072903, -0.016027, -0.009198, -0.007740, -0.008507, -0.021831, 0.021704, -0.001589, -0.002783, 0.003386, 0.008795, -0.053792, -0.069651, -0.064531, -0.099259, -0.159955, -0.177288, -0.085318, 0.031297, 0.120542, 0.168607, 0.044349, 0.022604, -0.056490, -0.053153, -0.071482, -0.087761, -0.052929, -0.083078, -0.069214, -0.049944, 0.020404, 0.012303, -0.026182, 0.017333, 0.032182, -0.036788, 0.021347, -0.009657, -0.028833, -0.018945, -0.045374, -0.094523, -0.106419, -0.130098, -0.087686, 0.016724, 0.230591, 0.234565, 0.132168, 0.001011, -0.065385, -0.123241, -0.130152, -0.061476, -0.044073, -0.021705, -0.034050, -0.014320, -0.010558, 0.024481, -0.015427, 0.022471, 0.024366, -0.033772, -0.002892, -0.018050, -0.046148, -0.030302, -0.077585, -0.079467, -0.167082, -0.152084, -0.146598, 0.063863, 0.329374, 0.361036, 0.129995, -0.069104, -0.084817, -0.126357, -0.086136, -0.087544, -0.046485, 0.003240, -0.043703, -0.037704, 0.005686, 0.004921, -0.006533, 0.031166, -0.021701, -0.022319, -0.028819, -0.017084, -0.031564, -0.019281, -0.073394, -0.103027, -0.181484, -0.173047, -0.112496, 0.090137, 0.398494, 0.300746, 0.072030, -0.113282, -0.133324, -0.066964, -0.100784, -0.013799, -0.022250, 0.014119, -0.025281, 0.021493, 0.003778, 0.002736, 0.024384, -0.033956, -0.028877, 0.034186, -0.023223, -0.035899, -0.024660, -0.055548, -0.078684, -0.149403, -0.176662, -0.258833, -0.148922, 0.207090, 0.427294, 0.284549, -0.009680, -0.151386, -0.147789, -0.111610, -0.083607, -0.056040, 0.010315, -0.022192, 0.003388, 0.022099, -0.003498, -0.019302, -0.024198, -0.013165, 0.012714, -0.030071, -0.005988, 0.002549, 0.003017, -0.037045, -0.071473, -0.107743, -0.179141, -0.213925, -0.111184, 0.221346, 0.382648, 0.206744, -0.097881, -0.196091, -0.137976, -0.078615, -0.080007, -0.075892, -0.047173, -0.035768, 0.010368, -0.026207, -0.003893, -0.007582, -0.021676, 0.016186, -0.014764, -0.002096, -0.027680, -0.017669, -0.026834, -0.053923, -0.095504, -0.119970, -0.189090, -0.180619, -0.027755, 0.277846, 0.328740, 0.151057, -0.177555, -0.222312, -0.153476, -0.101240, -0.077604, -0.024694, -0.054816, -0.008667, -0.011854, -0.033104, -0.014799, 0.008996, 0.006822, 0.025968, 0.024041, -0.020515, -0.019952, -0.026914, -0.068206, -0.074308, -0.119118, -0.108843, -0.103897, -0.070392, 0.044372, 0.266311, 0.295738, 0.045837, -0.175427, -0.197065, -0.125535, -0.095796, -0.069341, -0.058473, -0.018941, -0.010910, -0.046033, -0.027692, -0.000151, 0.013459, 0.017375, -0.021218, -0.035705, -0.003491, -0.011568, -0.018864, -0.069204, -0.052647, -0.091710, -0.071411, -0.082630, 0.018782, 0.132001, 0.253234, 0.238494, -0.041260, -0.130199, -0.182063, -0.148297, -0.090816, -0.071841, -0.037815, -0.015078, -0.054664, 0.006849, -0.013377, -0.009826, 0.007079, 0.027927, -0.019417, -0.024524, 0.019527, -0.028266, -0.028031, -0.082043, -0.083066, -0.059060, -0.075478, -0.025260, 0.072405, 0.140159, 0.193229, 0.106400, 0.010905, -0.133523, -0.161211, -0.146726, -0.103367, -0.051753, -0.053251, -0.009262, -0.030360, -0.021410, 0.014519, -0.001673, -0.007033, 0.011940, 0.028152, 0.008184, 0.021235, 0.008951, -0.035045, -0.065352, -0.077102, -0.063992, 0.007600, 0.051858, 0.073552, 0.080435, 0.138740, 0.041842, 0.010805, -0.073444, -0.096804, -0.106188, -0.104897, -0.035764, -0.062624, -0.025557, -0.001921, -0.044506, -0.001033, -0.013110, 0.025416, -0.022739, 0.021654, 0.021378, 0.015262, 0.020829, -0.030013, -0.084481, -0.028800, -0.026218, 0.008026, -0.003061, 0.021681, -0.007477, 0.050103, 0.046332, 0.013282, -0.028835, -0.097031, -0.089303, -0.078781, -0.067506, -0.012818, -0.017194, 0.011162, -0.010745, -0.034251, -0.010672, 0.025112, 0.021749, 0.011051, -0.011291, -0.035880, -0.025016, 0.012420, -0.019366, 0.015905, 0.026504, 0.013249, 0.037239, -0.042805, -0.066516, -0.064933, -0.040600, 0.014752, 0.000121, -0.050963, -0.024807, -0.080432, -0.074082, -0.051643, -0.036200, -0.018151, -0.012632, 0.015347, -0.031607, 0.005259, 0.000624, 0.009434, 0.034980, 0.020412, -0.019052, -0.008668, 0.024547, 0.027162, 0.064218, 0.038952, 0.016797, -0.066261, -0.119814, -0.077421, 0.005351, 0.036613, 0.063847, -0.016163, 0.001500, -0.050633, -0.055870, -0.028086, 0.001095, 0.016949, 0.006096, -0.003160, -0.001931, -0.014478, -0.003205, -0.002468, 0.030294, 0.019657, -0.025996, 0.021771, 0.021327, 0.049687, 0.026856, 0.042040, -0.049057, -0.044619, -0.061699, -0.079735, -0.029600, 0.053054, 0.040237, 0.034844, -0.032365, 0.000579, -0.043412, -0.029747, -0.025919, 0.013027, -0.002129, -0.034309, -0.020266, -0.016528, -0.033137, 0.004573, 0.012719, -0.007197, -0.015118, 0.004494, -0.020699, -0.022497, -0.017244, -0.005335, -0.080635, -0.074534, -0.107270, -0.088290, -0.088420, -0.003804, 0.010202, -0.015287, 0.011291, 0.021670, 0.011947, 0.015286, -0.036335, -0.034798, -0.027781, 0.011290, -0.030867, -0.027262, -0.017311, -0.032917, 0.000048, 0.005067, -0.021749, 0.020907, -0.019380, -0.024118, 0.004066, -0.003916, -0.052638, -0.077471, -0.067837, -0.045431, -0.022821, -0.018624, -0.039048, -0.046439, -0.037665, -0.015201, -0.001716, -0.017168, -0.028858, 0.003485, -0.028447, -0.027427, -0.029035, -0.009678, 0.031545, 0.013961, -0.004235, 0.007336, 0.013972, -0.000360, -0.030211, -0.024918, -0.028980, -0.007475, -0.041859, -0.017160, -0.024607, 0.021703, 0.017975, 0.013389, -0.003086, -0.014701, 0.007332, -0.025714, -0.015835, -0.007514, -0.008514, -0.033872, 0.014194, 0.029406, -0.019699, 0.009627, -0.004142, -0.001303, 0.002082, 0.030949, 0.004783, -0.022626, -0.012924, 0.017356, 0.011006, 0.000483, -0.005178, -0.014250, -0.013209, -0.019462, 0.005226, 0.009505, 0.026825, -0.008579, 0.002185, 0.022990, 0.015470, 0.004567, 0.010944, 0.001852, -0.030635, 0.001377, -0.007806, 0.032229
--  Sum of weights (converted): FFFFFFFE96129AAF
    );

    constant weights_n2 : weight_array := (
     x"01081546", x"003A0B1E", x"01058054", x"FF6951F6", x"00FE4B9E", x"00FBE651", x"FFF4D150", x"FF15356B", x"FFA19699", x"FFB1C227", x"0004D52B", x"FEF6BD60", x"00363ECC", x"FF8A321D", x"FFB95751", x"FF6910F6", x"FFC23A6E", x"FEF04814", x"FF64E354", x"001AF400", x"00BFB70C", x"0109DFA8", x"FF22AEC6", x"007ADB60", x"FF5B1426", x"FF1DCBDD", x"FFF31DD5", x"FF582AD9", x"FF04061F", x"FEEE94D2", x"FF3C2AF4", x"00F06A9A", x"00A3256F", x"FF8C1DBB", x"FF3B71B6", x"FF1CAE5D", x"FF51B2C8", x"FF82BEE3", x"00A7835D", x"00544DDF", x"FF83AAF0", x"00C60159", x"FF4DDC12", x"FF13FA43", x"004E7D4A", x"FF5E686A", x"004D7C6C", x"00F2B83B", x"FF71BB94", x"FF318BAD", x"006D597A", x"FEF79C0E", x"01050696", x"FF75D4D2", x"008D7250", x"FF175AFF", x"FF39F7BB", x"00203A64", x"0067FAD0", x"00E2C9D9", x"00F3D44A", x"FFEF0B97", x"FFD84BC7", x"002AD87D", x"FFB59905", x"000303F1", x"FED8FC4C", x"FEFE73CC", x"00B8B3C2", x"FF3AB306", x"00D0C246", x"00117CE5", x"002FBFF5", x"00D41E76", x"FF1006A3", x"FF7D05C0", x"FFF5F5D5", x"0035C9C5", x"FEC4EA08", x"005D660C", x"FF54B7A7", x"00291582", x"00C5F06A", x"FFE2DAFE", x"FFF6BE9C", x"FFEA23F3", x"00F42729", x"00A60B38", x"00302408", x"FF5650A7", x"FF716DD9", x"0122602E", x"014B9D72", x"019C266C", x"00779CBC", x"02948120", x"01CD3158", x"02DDB8C4", x"02BEFC20", x"019515D0", x"00AAD806", x"01955D9C", x"FF3D6012", x"0032EA15", x"FE4A8E4C", x"FF212C0C", x"FEA4ADE0", x"FF494709", x"006AB659", x"FF2DA1D8", x"FF027A9C", x"00D132EC", x"009C2E3E", x"FFFCC652", x"FF319659", x"FFB22AE2", x"FFA19395", x"00DE29AE", x"00166FF4", x"00A5C076", x"00ED8A55", x"02558C44", x"0462E188", x"0558C580", x"0560FB08", x"04D41780", x"06563C98", x"04FC5270", x"03BEC7B0", x"02605180", x"00F1F536", x"00476020", x"FF7BFDE4", x"FFAF6D24", x"FF06184A", x"005B8F4C", x"FF4540CF", x"FF6CB382", x"FF921FF9", x"FEED20E0", x"FF3FF1C4", x"FEF7426C", x"FFEEAEAB", x"00038B78", x"FFBC4F77", x"FF97702A", x"021BE848", x"01B69E18", x"03C0BB58", x"0534EBD0", x"0472C700", x"05731B48", x"06566DC0", x"06E38DA8", x"05C61698", x"06B64190", x"0483FDA8", x"0347ED1C", x"02E89CD4", x"00081398", x"0038AD53", x"FEDBF4BC", x"FE5D5292", x"000F447C", x"0078C096", x"FFF92DC4", x"FF49555E", x"FFF2CAEB", x"FF734C26", x"00D52E73", x"000D17AF", x"003EDF3C", x"00C922DB", x"00ED2EEE", x"00DD2296", x"03AB3C78", x"042FCFC8", x"033BD558", x"04CA41F8", x"03FDD70C", x"0346ACB4", x"02A1EBEC", x"03494C94", x"024AD518", x"03B99E90", x"031B52D4", x"00C8E79F", x"01084018", x"FEBF1C78", x"FF0315EA", x"FDEEB238", x"FE8E178E", x"FFB22566", x"003DAC2A", x"FFEC0BCB", x"FF6B6716", x"00CC80BC", x"00C0D16B", x"0033D102", x"FF799FA5", x"0066AD19", x"00BD0499", x"02EF1C20", x"028EBCE4", x"0290218C", x"022BDE04", x"02997C58", x"02004C94", x"02A30E44", x"0232F72C", x"00B32373", x"0124DA7E", x"FFED61AF", x"FF68F674", x"000DFE7C", x"FFCBDC83", x"FF22368F", x"0045D48E", x"FE630812", x"FDE67008", x"FEC51A80", x"FFA234D3", x"FFD831FF", x"01064BAA", x"FF845C86", x"FF67D466", x"001A54E5", x"00D61EC4", x"0078DD26", x"01731B36", x"01BE9748", x"02577BEC", x"018DE1C0", x"016F3A20", x"00FDC8F6", x"00214C84", x"00065D99", x"00BF396B", x"017ED23C", x"0052C37F", x"0179FDE2", x"00941779", x"FFF13460", x"FFCF1FAD", x"FF316346", x"004A4226", x"FEF23938", x"FF1FB9E7", x"FDCEA718", x"FEF13492", x"00103B59", x"00E8F5CD", x"008B1E90", x"0036C8A9", x"FEDE2214", x"0005A55C", x"FF72B43B", x"FFC14CE9", x"00B8490C", x"FEDB5952", x"FFA07F84", x"FE4BD9C0", x"FFCFCF43", x"FFC54D0E", x"FD8FE6C8", x"FEE60878", x"FEF77476", x"00CAB6F0", x"01FC3064", x"008A5769", x"0007BF9E", x"00C8F8E4", x"FFA9E040", x"FF1939D8", x"FFC4F6E3", x"FDE92918", x"FED2FCDA", x"0061BBA5", x"0063BEB5", x"FF419E82", x"004BC626", x"FF1FC2FB", x"FF5F46AB", x"00BF3424", x"FFAAB949", x"FF67C91C", x"FF4B1298", x"FDC74398", x"FBFECBF8", x"FBF8EDF8", x"FB818738", x"FC3710F0", x"FA7047A0", x"FB3A98D0", x"FC9248B0", x"FE066A28", x"FFFE8FAC", x"FFDC56C3", x"FFCFE8CC", x"FFF3D79C", x"FEB43908", x"FE4CBD4E", x"FFA989BC", x"FEBFC334", x"FEB82530", x"FFB5BFC5", x"00D01211", x"FF0B0605", x"FF64C407", x"FF2B7A07", x"FFE69EBF", x"FFE663CA", x"FEDBDB72", x"FFC6E9B4", x"FC64C8F4", x"FC816224", x"F9CAEF10", x"FA260D08", x"F9DC9978", x"F8432078", x"F9404320", x"F7F77850", x"FAA339B0", x"FC900994", x"FF76974A", x"003D04B4", x"009D7DD6", x"00433E30", x"FF1A41D5", x"00294DDC", x"FE83FCF2", x"FF4DD04E", x"FED2F072", x"FF67D8CA", x"FF0A1E14", x"010D0E2A", x"00307FED", x"FF2D6A00", x"0016B06A", x"FF611424", x"FF9323B3", x"FE7469D8", x"FB4E7770", x"FA5626A8", x"F8DD7ED8", x"F95A75F8", x"F752A680", x"F80468C0", x"F91620D8", x"F9E2D260", x"FAE14738", x"FD5E93AC", x"FEB4D260", x"FE5E985A", x"FF8BCD68", x"0042249A", x"008E4D12", x"FFA56D30", x"FD6C4368", x"FE138DBE", x"FED1C7C6", x"0086CC2B", x"FEFA0702", x"00693D74", x"FFAFB1FC", x"0069A694", x"0059EEA7", x"FF4F30F7", x"FFE953F1", x"FE063664", x"FA9677C0", x"FB7E9D18", x"FB3B7458", x"FAD7FDB0", x"F9EAB5B8", x"FAE93818", x"FA9B7E18", x"FB60C328", x"FCE8F330", x"FD3F4940", x"FDCC48B4", x"FD10C084", x"FFF1F9D4", x"FF01E78B", x"FFF8FEA1", x"FF254FCC", x"FE309C62", x"FF4C37E6", x"0014B620", x"00EF73DC", x"FFCFBFB9", x"011C8CD0", x"004CAC45", x"00AB3F6A", x"FFBC05AB", x"00B78E87", x"0070BC18", x"FCEBD438", x"FD875854", x"FB9C9C80", x"FC0C68D4", x"FC4A47C0", x"FE305D9A", x"FE0AA416", x"FF17A921", x"FF014224", x"FF3D1149", x"FD17E960", x"FE1432F8", x"FEA17998", x"FF4CFA39", x"FE678318", x"FF034645", x"FD491C98", x"FCF37A48", x"FE4AEA68", x"FEF60048", x"01212C88", x"FF844988", x"FFE99BE2", x"00798473", x"FEFD6DD0", x"00DE9746", x"FF7E1EDF", x"FF98BBEA", x"FE7B4E2C", x"FE55A880", x"FEA6111E", x"FEC405CA", x"00991ACF", x"00FCD4A4", x"030F5AD4", x"0357CFEC", x"0358D4FC", x"0127B98A", x"00B28433", x"01542C54", x"009D26DE", x"FE7A824A", x"FEDEB190", x"FD98AD00", x"FEA33A78", x"FE334D02", x"0034B259", x"0082C475", x"00E32E58", x"FF99B921", x"FF241074", x"002E0E23", x"FF6D2B1D", x"FF714AE4", x"0100921E", x"00116D82", x"00576D0C", x"0217F1E4", x"01B4CE22", x"00D779C8", x"028A4FC4", x"0385A1F0", x"02EFF15C", x"04E06028", x"04025CB8", x"0209A004", x"02F0E1CC", x"0161B3C2", x"01E2B5D4", x"FFADA8E4", x"FEF8FC8A", x"00A7A64F", x"FFC1F0F9", x"0078ABD1", x"017F13A0", x"008C2445", x"00A4FBAF", x"00F1AEBA", x"010C7B00", x"FFE10A93", x"00CD0F56", x"005ED87E", x"00C7151A", x"00D6C0E0", x"039B752C", x"03827AF4", x"02EF8A10", x"0377BFC4", x"02136B34", x"03DEC6C4", x"042F5E30", x"0507A9F0", x"04946018", x"0385FBA0", x"03432E60", x"01D6AD0E", x"01115216", x"011A723C", x"00BA3889", x"00679FD6", x"02EE6E50", x"0276DBC4", x"01E63EAA", x"036E0B58", x"02802784", x"FFE239F9", x"009A2CC7", x"FF4A7C70", x"0064F688", x"01005C5E", x"014A8FFE", x"02B11CB4", x"0362F410", x"044C6170", x"046A5500", x"03C7B874", x"038A57CC", x"04B1C850", x"049A1838", x"04C85650", x"03B0AD0C", x"02A0BD08", x"021234D0", x"039FE0C8", x"0230C050", x"009B2E09", x"01280574", x"0295FCE8", x"02C8A228", x"03809DCC", x"03EB0DB0", x"03724970", x"01E31652", x"004EC4CB", x"00C3FED3", x"00BB3807", x"00F00AC0", x"FFDCE390", x"FFED63A8", x"022FC184", x"02F01204", x"04ED13B8", x"047CACE8", x"04164038", x"03A9E834", x"0528F288", x"054BD570", x"053AD350", x"030D09DC", x"02A95C34", x"01D8DB64", x"00CE1ED9", x"00E2D2E2", x"02646CD4", x"01A071C4", x"03F25874", x"048B6630", x"051B8EE0", x"054589E8", x"03BF12E8", x"01E88574", x"00D5492B", x"FF87DCFA", x"FF64DAD4", x"FFC971C5", x"0091A68D", x"013BA1F6", x"02DAB938", x"02E4E9DC", x"0410BF28", x"03C952D4", x"05544678", x"03CEC5D8", x"034CA710", x"0407FD08", x"022F693C", x"00AA231D", x"FFD26491", x"FF99F8BE", x"019933E2", x"0043BD1D", x"036E6600", x"04663190", x"043AB4E0", x"04BDC048", x"05A5C760", x"046D3010", x"03922AF0", x"01BE6FAE", x"FF632F68", x"00B48373", x"00938AF9", x"FF3003DA", x"0083B98B", x"FFBB0100", x"00946117", x"023D1AB8", x"02DC06FC", x"0331C2FC", x"02E880CC", x"045782A8", x"03D71C9C", x"017BD202", x"FFD91B43", x"FF95DDFD", x"FDF9DD34", x"FE0AF586", x"FF909404", x"020BD034", x"01DEF34C", x"0395E3EC", x"03597A50", x"032701BC", x"0397F060", x"02E69A60", x"016D9604", x"014CD36A", x"0085AAB6", x"00B626C6", x"00729675", x"001EAF9F", x"009946AE", x"FF702EA9", x"013FE0C4", x"018C17F4", x"00E66C9E", x"01B5B3EA", x"010FF352", x"00CF688F", x"01191844", x"007402F7", x"FEFB9840", x"FE6D076E", x"FC969AC0", x"FD0F9730", x"FF9E04E1", x"FF1E4E5A", x"01EE25F0", x"0345AE8C", x"038EDF58", x"031EF724", x"01584396", x"01B27D86", x"004E4756", x"FFD9D2DD", x"00E05B6E", x"FF9C916E", x"FF2E7809", x"FF15244B", x"00B641B3", x"0006DBB5", x"011D4966", x"00285D6A", x"FE9EE1C0", x"FF81CC5D", x"FFB7B9DA", x"FEF10212", x"FE3EBBD0", x"FCB504B4", x"FC3A1B7C", x"FD043468", x"FB74C678", x"FCD2D1CC", x"FD585954", x"FEE35EE0", x"FFC08092", x"FF8C5DF6", x"0040C0BF", x"01EA8092", x"00E67910", x"0106081E", x"FF9BB178", x"00FA217B", x"FFC12492", x"FF9D6280", x"003B5974", x"FF972AF2", x"FF89740E", x"FFC39AC3", x"FFC340E3", x"FEF13508", x"FF8910A3", x"FD783FC8", x"FEA61EB4", x"FE7AF44E", x"FD532D24", x"FCE19278", x"FC302640", x"FDCF3C68", x"FE7097A0", x"FEB0078C", x"FE2E2608", x"FEEF1BB6", x"001330F0", x"FF63587D", x"FEF73EF2", x"FEB7B706", x"00708933", x"00726CD0", x"011CBDA2", x"FF7A33AF", x"007FABDE", x"FF9F3395", x"FFB74927", x"00AAB625", x"FEF3BE56", x"00D34C0A", x"00766C96", x"FF25C790", x"003BC905", x"FF102A12", x"FF25D6E0", x"FE9F008A", x"FDCCB074", x"FED17C62", x"FF886ED1", x"FEE563E6", x"FE91667C", x"FF46E63B", x"FF7C674F", x"FF09F90F", x"FE8B960E", x"FEE5271A", x"FF7A5187", x"002BC2D3", x"00DD6728", x"FFF2034C", x"006435E8", x"00AA1617", x"FF82907E", x"FF9EEB7B", x"00C2107A", x"00D17A4A", x"004553D0", x"FF1DD39B", x"00A3E1DC", x"FF08A5DB", x"0083B07B", x"0006F63E", x"00399612", x"FEBAA914", x"FF65B3B7", x"0040EFA7", x"00A5F5D3", x"FF723CCE", x"00D0A4D8", x"FF8FD5F3", x"FF21A546", x"FF59182D", x"FFF26BE5", x"FFB2EFB9", x"007AAFB6", x"FF540EFF", x"FFA9BC69", x"FEDD8F00", x"00EEBBE5", x"FFC8E26B", x"FF195CC6", x"FFF1E1DA", x"FFFF774A", x"0051415E", x"FFDFE317", x"00B80BC1", x"FF9B09D5", x"FFA82BE6", x"FFB9CC47", x"003368E6", x"00E96E74", x"FFF11C02", x"00DECF60", x"00E36D10", x"FF6442A8", x"FFE2CB3B", x"FF70CF28", x"007519FD", x"FF9484B1", x"0054A788", x"000ED959", x"FF3EF1D1", x"FF3A1768", x"FEE1BE78", x"FF5B9D5C", x"0051AFCC", x"0011D33D", x"00DC0B28", x"FEFEBCDA", x"FFF77357"
--  0.032237, 0.007085, 0.031922, -0.018394, 0.031042, 0.030749, -0.001365, -0.028661, -0.011525, -0.009551, 0.000590, -0.032380, 0.006622, -0.014380, -0.008625, -0.018425, -0.007540, -0.033169, -0.018935, 0.003290, 0.023403, 0.032455, -0.027016, 0.014997, -0.020132, -0.027613, -0.001573, -0.020487, -0.030759, -0.033376, -0.023905, 0.029348, 0.019915, -0.014146, -0.023994, -0.027749, -0.021277, -0.015290, 0.020448, 0.010291, -0.015177, 0.024171, -0.021746, -0.028811, 0.009581, -0.019726, 0.009459, 0.029629, -0.017367, -0.025202, 0.013348, -0.032274, 0.031863, -0.016866, 0.017266, -0.028399, -0.024174, 0.003934, 0.012693, 0.027684, 0.029764, -0.002070, -0.004847, 0.005230, -0.009082, 0.000368, -0.036013, -0.031439, 0.022547, -0.024085, 0.025483, 0.002135, 0.005829, 0.025893, -0.029294, -0.015988, -0.001226, 0.006566, -0.038463, 0.011401, -0.020909, 0.005015, 0.024162, -0.003558, -0.001130, -0.002668, 0.029804, 0.020269, 0.005877, -0.020713, -0.017404, 0.035446, 0.040480, 0.050311, 0.014601, 0.080628, 0.056298, 0.089566, 0.085814, 0.049449, 0.020855, 0.049483, -0.023758, 0.006215, -0.053399, -0.027201, -0.042398, -0.022305, 0.013026, -0.025680, -0.030947, 0.025537, 0.019065, -0.000394, -0.025197, -0.009501, -0.011526, 0.027119, 0.002739, 0.020233, 0.028997, 0.072943, 0.137070, 0.167086, 0.168088, 0.150890, 0.198027, 0.155801, 0.117039, 0.074258, 0.029536, 0.008713, -0.016114, -0.009836, -0.030506, 0.011177, -0.022796, -0.017981, -0.013412, -0.033554, -0.023444, -0.032317, -0.002114, 0.000433, -0.008263, -0.012764, 0.065907, 0.053542, 0.117277, 0.162710, 0.139011, 0.170301, 0.198050, 0.215278, 0.180431, 0.209748, 0.141112, 0.102530, 0.090895, 0.000986, 0.006919, -0.035650, -0.051108, 0.001864, 0.014740, -0.000833, -0.022298, -0.001612, -0.017176, 0.026023, 0.001598, 0.007675, 0.024553, 0.028953, 0.026994, 0.114653, 0.130836, 0.101054, 0.149690, 0.124736, 0.102377, 0.082266, 0.102698, 0.071635, 0.116409, 0.097085, 0.024525, 0.032257, -0.039171, -0.030873, -0.064612, -0.045155, -0.009504, 0.007528, -0.002436, -0.018139, 0.024964, 0.023537, 0.006325, -0.016403, 0.012534, 0.023073, 0.091688, 0.079924, 0.080094, 0.067855, 0.081236, 0.062537, 0.082404, 0.068721, 0.021867, 0.035749, -0.002273, -0.018437, 0.001708, -0.006365, -0.027074, 0.008524, -0.050411, -0.065620, -0.038440, -0.011449, -0.004859, 0.032019, -0.015093, -0.018575, 0.003214, 0.026138, 0.014754, 0.045301, 0.054515, 0.073179, 0.048570, 0.044828, 0.030980, 0.004065, 0.000777, 0.023343, 0.046731, 0.010103, 0.046142, 0.018078, -0.001806, -0.005966, -0.025221, 0.009065, -0.032932, -0.027377, -0.068524, -0.033056, 0.001981, 0.028438, 0.016982, 0.006687, -0.035384, 0.000689, -0.017248, -0.007654, 0.022496, -0.035724, -0.011658, -0.053241, -0.005883, -0.007165, -0.076184, -0.034420, -0.032293, 0.024745, 0.062035, 0.016887, 0.000946, 0.024533, -0.010513, -0.028171, -0.007206, -0.065288, -0.036745, 0.011930, 0.012176, -0.023240, 0.009250, -0.027373, -0.019620, 0.023340, -0.010410, -0.018581, -0.022086, -0.069426, -0.125147, -0.125863, -0.140438, -0.118278, -0.173794, -0.149097, -0.107143, -0.061717, -0.000176, -0.004353, -0.005870, -0.001484, -0.040500, -0.053132, -0.010554, -0.039091, -0.040021, -0.009064, 0.025399, -0.029904, -0.018949, -0.025943, -0.003098, -0.003126, -0.035662, -0.006969, -0.112697, -0.109206, -0.193978, -0.182855, -0.191821, -0.241806, -0.210905, -0.251041, -0.167575, -0.107417, -0.016774, 0.007449, 0.019225, 0.008208, -0.028045, 0.005042, -0.046388, -0.021751, -0.036751, -0.018573, -0.030015, 0.032844, 0.005920, -0.025706, 0.002770, -0.019400, -0.013289, -0.048289, -0.146672, -0.176984, -0.222962, -0.207707, -0.271161, -0.249462, -0.216049, -0.191062, -0.160000, -0.082205, -0.040427, -0.050953, -0.014184, 0.008074, 0.017371, -0.011056, -0.080534, -0.060113, -0.036892, 0.016455, -0.031979, 0.012847, -0.009803, 0.012897, 0.010978, -0.021583, -0.002768, -0.061742, -0.169132, -0.140794, -0.148992, -0.161134, -0.190099, -0.159031, -0.168519, -0.144438, -0.096564, -0.086025, -0.068813, -0.091705, -0.001712, -0.031018, -0.000855, -0.026695, -0.056566, -0.021946, 0.002528, 0.029230, -0.005890, 0.034735, 0.009359, 0.020904, -0.008298, 0.022407, 0.013762, -0.096212, -0.077228, -0.137132, -0.123485, -0.115933, -0.056596, -0.061201, -0.028362, -0.031096, -0.023795, -0.090831, -0.060034, -0.042789, -0.021853, -0.049864, -0.030850, -0.084825, -0.095279, -0.053355, -0.032471, 0.035300, -0.015102, -0.002733, 0.014834, -0.031564, 0.027172, -0.015854, -0.012606, -0.047448, -0.052044, -0.042228, -0.038571, 0.018690, 0.030863, 0.095624, 0.104469, 0.104594, 0.036099, 0.021792, 0.041525, 0.019184, -0.047545, -0.035316, -0.075113, -0.042575, -0.056238, 0.006433, 0.015963, 0.027732, -0.012485, -0.026848, 0.005622, -0.017924, -0.017420, 0.031320, 0.002127, 0.010672, 0.065423, 0.053321, 0.026303, 0.079384, 0.110063, 0.091790, 0.152390, 0.125288, 0.063675, 0.091905, 0.043177, 0.058925, -0.010051, -0.032106, 0.020465, -0.007576, 0.014730, 0.046762, 0.017107, 0.020140, 0.029502, 0.032773, -0.003779, 0.025032, 0.011578, 0.024302, 0.026215, 0.112727, 0.109678, 0.091741, 0.108368, 0.064870, 0.120944, 0.130782, 0.157186, 0.143112, 0.110105, 0.101951, 0.057456, 0.033364, 0.034478, 0.022732, 0.012649, 0.091605, 0.077009, 0.059356, 0.107183, 0.078144, -0.003634, 0.018820, -0.022157, 0.012325, 0.031294, 0.040352, 0.084120, 0.105829, 0.134324, 0.137980, 0.118130, 0.110638, 0.146702, 0.143810, 0.149455, 0.115317, 0.082121, 0.064722, 0.113266, 0.068451, 0.018943, 0.036135, 0.080809, 0.086991, 0.109450, 0.122443, 0.107701, 0.058971, 0.009615, 0.023925, 0.022854, 0.029302, -0.004286, -0.002272, 0.068330, 0.091805, 0.153940, 0.140219, 0.127716, 0.114491, 0.161248, 0.165507, 0.163431, 0.095342, 0.083174, 0.057722, 0.025161, 0.027688, 0.074759, 0.050835, 0.123333, 0.142017, 0.159614, 0.164739, 0.117074, 0.059634, 0.026036, -0.014665, -0.018939, -0.006660, 0.017780, 0.038529, 0.089200, 0.090444, 0.127044, 0.118326, 0.166538, 0.118991, 0.103107, 0.125975, 0.068287, 0.020769, -0.005567, -0.012455, 0.049951, 0.008269, 0.107226, 0.137475, 0.132166, 0.148163, 0.176487, 0.138329, 0.111593, 0.054497, -0.019142, 0.022035, 0.018011, -0.025389, 0.016080, -0.008422, 0.018113, 0.069959, 0.089359, 0.099824, 0.090882, 0.135682, 0.120009, 0.046365, -0.004748, -0.012956, -0.063249, -0.061162, -0.013601, 0.063942, 0.058466, 0.112047, 0.104673, 0.098512, 0.112297, 0.090650, 0.044627, 0.040628, 0.016317, 0.022235, 0.013988, 0.003746, 0.018710, -0.017556, 0.039048, 0.048351, 0.028128, 0.053431, 0.033197, 0.025318, 0.034313, 0.014162, -0.031788, -0.049191, -0.106616, -0.091847, -0.011961, -0.027551, 0.060321, 0.102256, 0.111190, 0.097530, 0.042024, 0.053038, 0.009556, -0.004660, 0.027387, -0.012138, -0.025578, -0.028669, 0.022248, 0.000837, 0.034825, 0.004927, -0.043105, -0.015405, -0.008823, -0.033080, -0.054842, -0.102903, -0.117907, -0.093237, -0.141995, -0.099265, -0.082965, -0.034745, -0.007751, -0.014115, 0.007904, 0.059876, 0.028134, 0.031986, -0.012244, 0.030534, -0.007673, -0.012038, 0.007245, -0.012797, -0.014471, -0.007372, -0.007415, -0.033056, -0.014518, -0.079071, -0.042222, -0.047491, -0.083597, -0.097464, -0.119122, -0.068453, -0.048756, -0.041012, -0.056867, -0.033312, 0.002343, -0.019123, -0.032319, -0.040074, 0.013737, 0.013968, 0.034758, -0.016333, 0.015585, -0.011816, -0.008876, 0.020839, -0.032746, 0.025793, 0.014456, -0.026638, 0.007298, -0.029277, -0.026631, -0.043091, -0.068764, -0.036928, -0.014596, -0.034498, -0.044751, -0.022595, -0.016064, -0.030033, -0.045461, -0.034527, -0.016319, 0.005342, 0.027027, -0.001707, 0.012233, 0.020762, -0.015312, -0.011851, 0.023689, 0.025571, 0.008463, -0.027609, 0.020005, -0.030194, 0.016075, 0.000850, 0.007030, -0.039714, -0.018835, 0.007927, 0.020259, -0.017305, 0.025469, -0.013692, -0.027143, -0.020374, -0.001658, -0.009407, 0.014976, -0.020989, -0.010530, -0.035454, 0.029142, -0.006728, -0.028154, -0.001723, -0.000065, 0.009919, -0.003920, 0.022467, -0.012324, -0.010721, -0.008570, 0.006276, 0.028495, -0.001818, 0.027198, 0.027762, -0.019011, -0.003565, -0.017479, 0.014295, -0.013120, 0.010334, 0.001813, -0.023566, -0.024159, -0.034943, -0.020067, 0.009972, 0.002176, 0.026861, -0.031404, -0.001044
--  Sum of weights (converted): 00000000B2284934
    );

    constant weights_n3 : weight_array := (
     x"FEF9AA76", x"0001B66D", x"006A9830", x"FEF98CFC", x"0102629C", x"FFA52145", x"01033A98", x"FFCEE43E", x"00A5FAEA", x"0109F848", x"FF957B85", x"FFB8E139", x"009968E4", x"FF0521F9", x"00ACE0B9", x"FF483828", x"010FBACA", x"FF404242", x"FF879A80", x"00DA5003", x"FF809E47", x"00FAC72A", x"00C94B7C", x"010B69E6", x"FEE46A70", x"00034772", x"FF9FC4F0", x"0045B10B", x"FF2317F6", x"0077F857", x"FFF223CA", x"FF75B46D", x"FEF8CD04", x"0099084B", x"FF95F7AC", x"00D76C10", x"0033512C", x"00581284", x"FFD2FB7A", x"FFD6464C", x"FF9AB8A8", x"FF00AC6E", x"00B5F194", x"FF45E4F7", x"00A8AB43", x"FF9BEC31", x"00B69D8A", x"00FA5B3C", x"FF4CACB6", x"00F16AAF", x"000718DA", x"FF207DEF", x"00776E5C", x"00A5AA5A", x"0101E7B8", x"FEE97ECC", x"01082E56", x"00DDCCEE", x"011FD208", x"009F69EA", x"FF719F65", x"00DDE50E", x"010AEDB2", x"FF8E449B", x"FFCBF32B", x"00DD01BA", x"00E0F9FA", x"00B8146D", x"00D2E151", x"FF54DF25", x"FFB5B4EA", x"FF6FE9F2", x"007FCB80", x"00330EDF", x"FF080E81", x"FFC6FE9F", x"FF0375AD", x"FEE37A76", x"0105346C", x"FF6AD5CF", x"00820CF8", x"FFBED146", x"FFC4C127", x"FFFFCFA0", x"00E42F3E", x"FFD786DE", x"00F21690", x"00AB0B30", x"00C83ED6", x"FF017A66", x"FF806E84", x"FF1F7105", x"FFD5FA37", x"FFDD8D7E", x"006C60C1", x"0182D12A", x"0148407A", x"00061DEC", x"0032DE7D", x"01A253C2", x"00A86D1C", x"00B6CC2C", x"FF9D1866", x"FFDAC009", x"003E3B6B", x"FF107B83", x"0098F6CC", x"007D6C25", x"FF4C4EEC", x"FF86DBBB", x"FFBB0034", x"002D8822", x"FF94ADD0", x"0117EDCE", x"FEE65BF6", x"FF5D1D5B", x"FF5F65D2", x"00947173", x"00AE1DF9", x"00916ADB", x"02645320", x"00E87030", x"02DA07D4", x"02353CC4", x"028E271C", x"0172DDA8", x"00FC5067", x"00220F9E", x"00D1AD19", x"FF4BB90F", x"002EFD6B", x"FE997EE4", x"FEA2C980", x"FF0B294C", x"0022EE9D", x"FF14803C", x"00701995", x"00472E10", x"00B04CF6", x"00B8BFD7", x"0076BAEC", x"FFA7C6A0", x"FFAEDAB7", x"0085D847", x"00FF5E57", x"00ED8907", x"024CC454", x"01D44766", x"03F05FF0", x"03C25C9C", x"0383AE5C", x"03AA4120", x"02E5F954", x"036DA374", x"01C1B08C", x"01A61D32", x"01154224", x"FF11EDAA", x"FF411010", x"FECF0360", x"FEF0115E", x"FEF0D8E6", x"FD7FD374", x"FF47BBC5", x"FF5CF597", x"FF34A315", x"FF75CF06", x"004A4B4C", x"003CEAD4", x"FFF6A251", x"FF7174AD", x"00D8DB63", x"01178AF0", x"00AE6AD8", x"0292AA9C", x"031E3B58", x"03BC36D8", x"041CB2C0", x"03C1BC78", x"054AE3B8", x"02BAF558", x"04ADE400", x"02A659D8", x"0328A500", x"025B0C94", x"00F1584D", x"015021EC", x"00E7FBDD", x"FF50C2D9", x"FE8A224A", x"FEC0C9DC", x"FE141888", x"FF4BA9ED", x"00488A60", x"FF8742B3", x"FF5C7802", x"006BB175", x"FF98A137", x"FF3F359B", x"FFD3179B", x"00D6EE81", x"0368FDD0", x"0317FB3C", x"036985F0", x"03141A8C", x"01F1461E", x"02EEB6C0", x"0197A194", x"017DE580", x"02DBDCDC", x"023A630C", x"03C57434", x"02270000", x"02C62B54", x"01CDD4B2", x"00A3EFD8", x"022C6434", x"004F00A5", x"FE1EAE0C", x"FF133033", x"FF33E7B5", x"FFF37FB6", x"FF827251", x"FF5E934D", x"FF629163", x"006C8165", x"004703EC", x"FFB55F3A", x"026EE390", x"02A17664", x"018F9544", x"01F5CCA8", x"FFF4507B", x"FFEE8710", x"FFD3577A", x"FD54AB04", x"FDF92BE0", x"FF608E2C", x"016CCD06", x"01FCE03A", x"0269BDDC", x"022A2F9C", x"01B1A442", x"026ECE4C", x"027AE6BC", x"01328E92", x"FF75A746", x"FE4BDCE6", x"FEA73F56", x"FFF15311", x"00B71D67", x"FF6DB4D7", x"FF68143B", x"007D9575", x"FF2498B1", x"010A2D74", x"01717B60", x"012194B4", x"000CCFBD", x"FF5561CD", x"FCBE7530", x"FB1633C0", x"FBF28808", x"F9431110", x"FA5A7AF8", x"FD363488", x"00E6A621", x"03A1ECB0", x"03355DE8", x"02A415F4", x"01EC3972", x"0349D6E4", x"035B9190", x"016B4E96", x"FF8D163B", x"FF86E343", x"FE2894CE", x"002FF9C3", x"FF4AF705", x"00E39F91", x"FEFCD232", x"0068105C", x"FF0544EA", x"00E6D5E5", x"0083912C", x"00D918E6", x"FDF35E30", x"FDBCBC5C", x"FA4517B0", x"F8B59B68", x"F895A8F8", x"F853AA48", x"FA1A7AF0", x"FE3B9C22", x"0277FF78", x"04EE40B8", x"05914BE0", x"044D7768", x"02B81A44", x"01906CD2", x"009401FD", x"012C688A", x"FE8D1BA2", x"FEDB4D9A", x"FE905BE8", x"FF12A113", x"00321DEE", x"FFB77FA7", x"00212DFB", x"FFF8CDC7", x"0003BA74", x"FFDF13F5", x"FFE8F726", x"FF9463FB", x"FE77178C", x"FC8CC42C", x"F8F0D590", x"F816B0D0", x"F8E4F390", x"FAC452A0", x"FEF09936", x"03233894", x"04E62AE8", x"04A26200", x"04976898", x"046214E8", x"02E49F5C", x"0095E6C9", x"001FDA2A", x"FDAD1ECC", x"FE397462", x"FFEA79B2", x"FF23005E", x"00A5C189", x"FF0E1545", x"01029C1C", x"008B79D2", x"00BA1AB3", x"0041F514", x"0003D896", x"FF2C2F36", x"FE323ADE", x"FC897958", x"FC99E124", x"FA4AD8F0", x"FAFE4198", x"FB3544E0", x"FEED9970", x"0197A1E6", x"03861E88", x"05BFCD80", x"041BC350", x"0443F8D0", x"02063360", x"021A3660", x"FEC685C8", x"FE98330C", x"FE7DF4B2", x"FD889364", x"FFD20ED2", x"00995241", x"FF47BCB4", x"001727DC", x"00587A44", x"00F24B1F", x"00E286C3", x"FF02D4C6", x"FF05C8C2", x"FEB0B7BC", x"FE5D2A14", x"FD6A312C", x"FBED6918", x"FCC16440", x"FBC43330", x"FD1FC840", x"000D62DA", x"035D1DC4", x"0606F3D8", x"0456FA08", x"02F66BD4", x"02F7BF08", x"01AAA3FC", x"00AA6A27", x"FFBAFDCE", x"FF140165", x"FF1AEAC2", x"FE91ABD8", x"FE6C6618", x"FEF05CEE", x"0111F55A", x"FEF62B5C", x"00448594", x"FFE3BBBF", x"011151CA", x"00A92687", x"FFB5ACC3", x"FEDF7FDE", x"FF3A6F5D", x"FD1B0008", x"FCC9A4D8", x"FCFFC4F4", x"FDAAFFA8", x"FE196D44", x"002BA5FD", x"025818E8", x"01B81DB2", x"01E994DE", x"007F6740", x"01B7A15C", x"0192B7E4", x"00FFEB81", x"0145CB00", x"0074DEED", x"0058B9C7", x"00231522", x"FE552A8E", x"FEF642E4", x"FF0F1A32", x"00BFFB97", x"00ABF1B2", x"00ECF455", x"FF37E024", x"FF6DE7FB", x"013A37C0", x"FF318D04", x"FEB2147A", x"FEC935DA", x"FC415870", x"FC18CABC", x"FCD003B4", x"FE3D82C8", x"FF3233C0", x"FF8384C7", x"008F1802", x"00250B31", x"FE45F178", x"000D25A1", x"00A9AC1E", x"01CD4DA6", x"029FB5DC", x"02692E18", x"01790F74", x"FF065333", x"FF406647", x"0019DB9A", x"FFC3C640", x"FFA0D2B2", x"FF684BB0", x"011561B2", x"FF19D1B9", x"FF3F259D", x"0141EF36", x"FFEA49DF", x"00A399D5", x"FE1ADB26", x"FD66EBF4", x"FB96D1F0", x"FC3A8620", x"FBEB5550", x"FC1DA744", x"FCAB0964", x"FBE76E88", x"FB507478", x"FC75F608", x"FF8CE4B2", x"015DC8F8", x"03E82598", x"035EFD64", x"02BCAF30", x"01770788", x"0156A022", x"FED3F758", x"FFE9B604", x"003A629F", x"002C2759", x"00CD05E9", x"00463815", x"FFB15B5F", x"FF68EE31", x"FFD0BE15", x"01E089F8", x"012C37C6", x"FE561AC2", x"FE38EF88", x"FBCBA860", x"FB417068", x"F8FA2EA0", x"FA4F5ED0", x"FA8488D0", x"FA3380C0", x"FA8C6928", x"FC849C14", x"0002C349", x"0192FB24", x"032CB3E4", x"0380CFD8", x"036745C8", x"02219AD4", x"01E15C1A", x"00D1DED1", x"FFE7868D", x"0054DF19", x"FFD109EA", x"008B9A88", x"FF9B6988", x"00FED8F6", x"00472A9E", x"016BF8B4", x"0145E890", x"02D69EF4", x"0037DDCC", x"FF9E73A2", x"FC457BF8", x"F9E8BF68", x"F973FBC8", x"F88CC208", x"F992A2F0", x"F95D6A50", x"F99A6960", x"FDE1A4B8", x"01C51564", x"023BB880", x"031E404C", x"04638520", x"0264BDF4", x"02F6A514", x"0110E944", x"FFFD1D98", x"FEA56E40", x"FFC2B330", x"FF908221", x"FF7BD690", x"FF702828", x"00433155", x"0123A7BE", x"01ED20E0", x"03076ED4", x"041037B8", x"02C5EDDC", x"00578684", x"FDE6ED88", x"FD220D40", x"FC00B65C", x"FA2AF6B0", x"F9F540C0", x"FB814DC0", x"FDA2B1E8", x"FE035082", x"0153E79C", x"03579EE4", x"0318AAD4", x"031274CC", x"03F9F148", x"03303B3C", x"FFE0FC92", x"FF7F8E75", x"FE75DDFE", x"0045D8C3", x"FF30A5D6", x"FF6AB259", x"FF7863D6", x"002D077B", x"01242446", x"0193F700", x"03A9A16C", x"04DF3788", x"03333070", x"0250F4D0", x"013BCFFC", x"FF92331A", x"FEB39B76", x"FDEA9A5C", x"FC8747E0", x"FED59BB6", x"FFDAE9D2", x"00A30BE1", x"037D289C", x"0383FDBC", x"0467CC90", x"022D5A34", x"03A7D84C", x"025F5FA4", x"FEFA3A70", x"FE47635E", x"FF286133", x"FF2A88E7", x"0049ED8D", x"008236E1", x"FFDAB675", x"00CF059E", x"006294D7", x"013ADA48", x"020291F4", x"043D10C0", x"030C7E24", x"03890B18", x"02F7801C", x"00BC26FC", x"00710788", x"FF408850", x"FFC60EA2", x"006D7696", x"FFD864FB", x"010C8C10", x"023E4A5C", x"01E8A148", x"030D7AA4", x"017C821E", x"00612190", x"0043DEFC", x"FFF269FA", x"FEF525AA", x"FE78B8F0", x"00130E36", x"00938E28", x"00E48C33", x"001BC047", x"00CB2FE5", x"FF371669", x"0216020C", x"016D49C0", x"0235F830", x"04A27E18", x"039B66F0", x"0414D0A8", x"0248A7C4", x"03249098", x"02AF3E60", x"01743476", x"0245F384", x"00BC7FB5", x"0181AF70", x"01DD27B4", x"01FB2A20", x"008A2956", x"0184E874", x"FF961B42", x"FEB83BAC", x"FF98125B", x"FEADBA12", x"FEC3C678", x"005690EA", x"00636EE3", x"007081A9", x"FFD9A1F3", x"FF2A083B", x"FF2BD03D", x"019F69A0", x"006C4870", x"02986FE8", x"04108660", x"047F2D60", x"02C2128C", x"033437F8", x"0267A01C", x"0395B770", x"0139DD10", x"011A412C", x"0094AC19", x"01997EAA", x"00B2913E", x"00DB961B", x"0124C674", x"FF5654B3", x"FED0125E", x"FEBE2422", x"FFFA5522", x"003D75AD", x"002CC262", x"FF1A8984", x"001A42FA", x"FF64BFE9", x"FFC67779", x"FFD2B510", x"00136823", x"FF357436", x"01A0AC3A", x"00AF9E55", x"0238E320", x"03402C88", x"034C9E9C", x"03E15FF8", x"03DF9898", x"03E5F138", x"02DA3B08", x"03078ABC", x"00D73BBB", x"FFE7D32F", x"00A753FF", x"00109CEA", x"FF6407E0", x"FE859C4E", x"FFF3F0D0", x"007AF95C", x"FFB76EE7", x"0030201C", x"00797C89", x"FEDD0FA8", x"FFCFD4FD", x"FF93775B", x"FF6A761B", x"00B2D275", x"01228A12", x"002FC76B", x"00CAC888", x"FF576E6F", x"008CE141", x"005C6B83", x"00143859", x"012FDC00", x"0179C9D2", x"011EE18C", x"01B90A52", x"0183D73C", x"01865C86", x"001794DE", x"FFCAE20E", x"FF89DE8F", x"FFCDC919", x"FF174CDA", x"FFB75966", x"FEF04624", x"FF287392", x"FF012E44", x"00D77DD2", x"FF57C704", x"FFE861FF", x"001F4749", x"0102676A", x"0084C7D5", x"FF2FA672", x"011E1E00", x"FEEA3D78", x"00266FEE", x"01090414", x"00F987F7", x"FFAA6752", x"FF1DEDCA", x"004E6AD2", x"00A2F622", x"FF1F6F0B", x"FF8990DF", x"FEF6AA2C", x"00185D25", x"FFEF6018", x"00505775", x"FF756AEE", x"FED3EB80", x"FF7C6F74", x"FF169587", x"FFB861FD", x"0069E77B", x"FF0C8631", x"FFF25469", x"FEE1C100", x"FF30AB5F", x"FF3328CF", x"FF9C623B", x"FF6BC2B2", x"002D08A9", x"00B2D842", x"00DC6322", x"005BA22A", x"FFFD659A", x"FFCA93D9", x"00C45889", x"FF548C4A", x"00CF42BC", x"FEDFCB8C", x"FF1BCA37", x"003F6CE9", x"FF79C9C7", x"00266350", x"00F032F7", x"007C70EE", x"011A17EE", x"FF8250B6", x"FF73A033", x"FFDA6289", x"FFC50880", x"FF7F4E82", x"FFEDD5DA", x"0108509C", x"FF5F9FED"
--  -0.032023, 0.000209, 0.013012, -0.032037, 0.031541, -0.011093, 0.031644, -0.005995, 0.020261, 0.032467, -0.013003, -0.008682, 0.018727, -0.030623, 0.021103, -0.022434, 0.033170, -0.023406, -0.014697, 0.026649, -0.015550, 0.030613, 0.024572, 0.032643, -0.034617, 0.000400, -0.011747, 0.008507, -0.026966, 0.014645, -0.001692, -0.016882, -0.032129, 0.018681, -0.012943, 0.026297, 0.006264, 0.010751, -0.005495, -0.005093, -0.012363, -0.031168, 0.022210, -0.022718, 0.020589, -0.012216, 0.022292, 0.030561, -0.021890, 0.029470, 0.000866, -0.027284, 0.014579, 0.020223, 0.031483, -0.033997, 0.032249, 0.027075, 0.035134, 0.019460, -0.017380, 0.027087, 0.032584, -0.013883, -0.006354, 0.026978, 0.027463, 0.022471, 0.025742, -0.020890, -0.009069, -0.017589, 0.015600, 0.006233, -0.030267, -0.006959, -0.030828, -0.034732, 0.031885, -0.018209, 0.015875, -0.007957, -0.007232, -0.000023, 0.027855, -0.004941, 0.029552, 0.020879, 0.024444, -0.031070, -0.015572, -0.027412, -0.005130, -0.004205, 0.013230, 0.047219, 0.040070, 0.000747, 0.006210, 0.051065, 0.020560, 0.022314, -0.012073, -0.004547, 0.007597, -0.029238, 0.018672, 0.015310, -0.021935, -0.014788, -0.008423, 0.005558, -0.013101, 0.034171, -0.034380, -0.019883, -0.019605, 0.018121, 0.021255, 0.017751, 0.074747, 0.028374, 0.089115, 0.068999, 0.079853, 0.045272, 0.030800, 0.004158, 0.025595, -0.022006, 0.005736, -0.043763, -0.042629, -0.029888, 0.004264, -0.028747, 0.013684, 0.008689, 0.021521, 0.022552, 0.014493, -0.010770, -0.009905, 0.016338, 0.031173, 0.028996, 0.071871, 0.057163, 0.123093, 0.117476, 0.109824, 0.114533, 0.090573, 0.107134, 0.054894, 0.051528, 0.033845, -0.029061, -0.023308, -0.037230, -0.033195, -0.033100, -0.078146, -0.022493, -0.019902, -0.024825, -0.016869, 0.009069, 0.007436, -0.001143, -0.017400, 0.026472, 0.034124, 0.021291, 0.080404, 0.097440, 0.116725, 0.128503, 0.117399, 0.165392, 0.085322, 0.146227, 0.082807, 0.098711, 0.073614, 0.029461, 0.041032, 0.028318, -0.021391, -0.045638, -0.038966, -0.060047, -0.022014, 0.008855, -0.014739, -0.019962, 0.013146, -0.012618, -0.023534, -0.005482, 0.026237, 0.106566, 0.096677, 0.106631, 0.096204, 0.060702, 0.091640, 0.049760, 0.046618, 0.089339, 0.069627, 0.117853, 0.067261, 0.086691, 0.056376, 0.020012, 0.067919, 0.009644, -0.058755, -0.028908, -0.024914, -0.001526, -0.015326, -0.019705, -0.019218, 0.013245, 0.008669, -0.009110, 0.076036, 0.082210, 0.048777, 0.061255, -0.001426, -0.002133, -0.005451, -0.083415, -0.063334, -0.019463, 0.044531, 0.062119, 0.075408, 0.067650, 0.052935, 0.076026, 0.077503, 0.037421, -0.016888, -0.053239, -0.042084, -0.001791, 0.022353, -0.017858, -0.018545, 0.015330, -0.026783, 0.032492, 0.045103, 0.035349, 0.001564, -0.020827, -0.101751, -0.153540, -0.126644, -0.210563, -0.176455, -0.087133, 0.028155, 0.113516, 0.100265, 0.082530, 0.060086, 0.102764, 0.104928, 0.044349, -0.014027, -0.014784, -0.057546, 0.005856, -0.022099, 0.027786, -0.031638, 0.012703, -0.030607, 0.028178, 0.016060, 0.026501, -0.064042, -0.070711, -0.179066, -0.227831, -0.231731, -0.239787, -0.184268, -0.055223, 0.077148, 0.154084, 0.173986, 0.134456, 0.084973, 0.048880, 0.018067, 0.036671, -0.045275, -0.035730, -0.044878, -0.028976, 0.006118, -0.008850, 0.004050, -0.000878, 0.000455, -0.004019, -0.002812, -0.013136, -0.047962, -0.107817, -0.220601, -0.247230, -0.222052, -0.163535, -0.033130, 0.098049, 0.153097, 0.144822, 0.143482, 0.136973, 0.090408, 0.018299, 0.003888, -0.072617, -0.055486, -0.002628, -0.026977, 0.020234, -0.029531, 0.031569, 0.017026, 0.022718, 0.008051, 0.000469, -0.025856, -0.056368, -0.108219, -0.106216, -0.178363, -0.156463, -0.149747, -0.033496, 0.049760, 0.110122, 0.179663, 0.128389, 0.133297, 0.063257, 0.065700, -0.038266, -0.043921, -0.047125, -0.077078, -0.005608, 0.018716, -0.022493, 0.002827, 0.010800, 0.029577, 0.027652, -0.030904, -0.030544, -0.040928, -0.051127, -0.080787, -0.127269, -0.101393, -0.132300, -0.089870, 0.001634, 0.105117, 0.188349, 0.135617, 0.092581, 0.092742, 0.052080, 0.020803, -0.008424, -0.028808, -0.027964, -0.044718, -0.049268, -0.033159, 0.033442, -0.032450, 0.008364, -0.003451, 0.033364, 0.020648, -0.009073, -0.035217, -0.024117, -0.090454, -0.100385, -0.093778, -0.072876, -0.059396, 0.005328, 0.073254, 0.053725, 0.059763, 0.015552, 0.053666, 0.049160, 0.031240, 0.039770, 0.014266, 0.010831, 0.004283, -0.052104, -0.032439, -0.029406, 0.023435, 0.020989, 0.028925, -0.024429, -0.017834, 0.038357, -0.025201, -0.040762, -0.037938, -0.117023, -0.121974, -0.099608, -0.054991, -0.025122, -0.015195, 0.017468, 0.004522, -0.053962, 0.001605, 0.020712, 0.056311, 0.081996, 0.075339, 0.046028, -0.030478, -0.023389, 0.003156, -0.007352, -0.011618, -0.018519, 0.033860, -0.028098, -0.023542, 0.039299, -0.002650, 0.019971, -0.059222, -0.081186, -0.137839, -0.117856, -0.127523, -0.121380, -0.104121, -0.127999, -0.146429, -0.110600, -0.014051, 0.042698, 0.122088, 0.105345, 0.085533, 0.045780, 0.041824, -0.036625, -0.002721, 0.007127, 0.005390, 0.025027, 0.008572, -0.009600, -0.018441, -0.005769, 0.058660, 0.036648, -0.051989, -0.055550, -0.131389, -0.148262, -0.219460, -0.177811, -0.171321, -0.181213, -0.170360, -0.108812, 0.000337, 0.049192, 0.099207, 0.109474, 0.106357, 0.066602, 0.058760, 0.025619, -0.002988, 0.010360, -0.005733, 0.017041, -0.012279, 0.031109, 0.008687, 0.044430, 0.039784, 0.088699, 0.006820, -0.011908, -0.116518, -0.190338, -0.204592, -0.232818, -0.200850, -0.207347, -0.199901, -0.066206, 0.055308, 0.069790, 0.097443, 0.137148, 0.074798, 0.092608, 0.033314, -0.000352, -0.042306, -0.007483, -0.013610, -0.016133, -0.017559, 0.008202, 0.035602, 0.060196, 0.094657, 0.126980, 0.086661, 0.010684, -0.065561, -0.089593, -0.124913, -0.182255, -0.188812, -0.140466, -0.073890, -0.062095, 0.041492, 0.104446, 0.096761, 0.096003, 0.124261, 0.099638, -0.003786, -0.015679, -0.048112, 0.008526, -0.025312, -0.018226, -0.016554, 0.005497, 0.035662, 0.049312, 0.114457, 0.152248, 0.099999, 0.072382, 0.038551, -0.013403, -0.040575, -0.065112, -0.108486, -0.036425, -0.004527, 0.019903, 0.109028, 0.109862, 0.137671, 0.068036, 0.114239, 0.074142, -0.031955, -0.053786, -0.026321, -0.026058, 0.009024, 0.015895, -0.004552, 0.025271, 0.012034, 0.038434, 0.062814, 0.132454, 0.095275, 0.110479, 0.092712, 0.022968, 0.013798, -0.023373, -0.007073, 0.013362, -0.004835, 0.032782, 0.070104, 0.059647, 0.095395, 0.046449, 0.011857, 0.008285, -0.001658, -0.032575, -0.047763, 0.002326, 0.018012, 0.027899, 0.003388, 0.024803, -0.024525, 0.065187, 0.044591, 0.069088, 0.144836, 0.112720, 0.127541, 0.071369, 0.098213, 0.083892, 0.045435, 0.071039, 0.023010, 0.047081, 0.058246, 0.061910, 0.016865, 0.047474, -0.012926, -0.040011, -0.012687, -0.041293, -0.038602, 0.010567, 0.012138, 0.013734, -0.004684, -0.026119, -0.025902, 0.050710, 0.013218, 0.081108, 0.127017, 0.140525, 0.086190, 0.100124, 0.075150, 0.112026, 0.038313, 0.034455, 0.018148, 0.049987, 0.021798, 0.026805, 0.035739, -0.020712, -0.037101, -0.039289, -0.000692, 0.007502, 0.005464, -0.028011, 0.003206, -0.018951, -0.007023, -0.005529, 0.002369, -0.024725, 0.050863, 0.021438, 0.069444, 0.101584, 0.103103, 0.121262, 0.121044, 0.121819, 0.089139, 0.094671, 0.026274, -0.002951, 0.020426, 0.002028, -0.019039, -0.046190, -0.001472, 0.015011, -0.008858, 0.005875, 0.014830, -0.035515, -0.005880, -0.013249, -0.018254, 0.021829, 0.035466, 0.005832, 0.024754, -0.020577, 0.017197, 0.011282, 0.002468, 0.037092, 0.046117, 0.035020, 0.053838, 0.047344, 0.047652, 0.002879, -0.006484, -0.014420, -0.006130, -0.028406, -0.008869, -0.033170, -0.026312, -0.031106, 0.026305, -0.020535, -0.002883, 0.003818, 0.031543, 0.016209, -0.025433, 0.034926, -0.033906, 0.004692, 0.032351, 0.030460, -0.010449, -0.027597, 0.009572, 0.019893, -0.027413, -0.014457, -0.032390, 0.002974, -0.002029, 0.009807, -0.016917, -0.036631, -0.016060, -0.028493, -0.008742, 0.012928, -0.029721, -0.001669, -0.034942, -0.025309, -0.025005, -0.012160, -0.018096, 0.005497, 0.021832, 0.026903, 0.011186, -0.000318, -0.006521, 0.023968, -0.020929, 0.025300, -0.035181, -0.027858, 0.007742, -0.016383, 0.004686, 0.029321, 0.015191, 0.034435, -0.015342, -0.017136, -0.004592, -0.007198, -0.015710, -0.002217, 0.032265, -0.019577
--  Sum of weights (converted): 00000000856AE45C
    );

    constant weights_n4 : weight_array := (
     x"00A44D9A", x"0087E9AE", x"00A96EF0", x"004EEE27", x"FF93EB72", x"0078BF89", x"FF76333B", x"FF4C6A24", x"01117E8C", x"00F28243", x"FF2C8EC2", x"00EDA465", x"003BC2EF", x"0048327E", x"0119187C", x"FFF0999B", x"FFA2F2BB", x"00B7AB53", x"FFB46CBB", x"FFB9C3CB", x"FF8A04E0", x"011FF98C", x"008B9A83", x"FFD09229", x"FFFA29C0", x"001479F6", x"FF52908F", x"00531177", x"FF1CED4F", x"FFF25BDC", x"FFC91A77", x"FF8889CB", x"010E91F8", x"0051D221", x"0089BA6F", x"FF381B03", x"00243D76", x"0043A248", x"0083EAF0", x"FF8DD911", x"FFA3F7D8", x"FEFA96AA", x"00A36181", x"00B2B135", x"00764706", x"008932D8", x"00A87407", x"010F0406", x"005BCB14", x"00666C0D", x"0059A87C", x"FF59BF58", x"004967D0", x"0058263E", x"FF17207F", x"FFA96969", x"FF4B7C2B", x"FF450F0F", x"00CB5140", x"00E61395", x"FFD68324", x"00593B0B", x"FFB662E0", x"0027F128", x"FFA96B83", x"FF2CBB4E", x"FF1C4C83", x"00904907", x"FF7D7EDC", x"FEB45C04", x"FF82CD51", x"FE4AC48E", x"FF835A11", x"007D18BC", x"FFD7FF8C", x"001B3CD0", x"FED309D2", x"FFB3F301", x"009EC996", x"FF231038", x"FF7444AE", x"00C4AC9E", x"00540530", x"0088C4F5", x"FEEF2C12", x"00BA34F7", x"FFC02CC8", x"003D04E1", x"00EBAF3B", x"FEEFC5B4", x"0046BFB8", x"FED12B1A", x"00887343", x"FFC6E234", x"FF40B78B", x"FE5ABB34", x"FEFA3DF2", x"FDCE2120", x"FE9E93A4", x"FF68D399", x"FDC64AE4", x"FE86F610", x"FF6C10AC", x"FFAE7ACC", x"FFBEE6D0", x"00D4352C", x"FF9D3380", x"0045B2A6", x"009478EC", x"FFC5A2C0", x"00BEE67E", x"00BF140E", x"0082482E", x"FFB89E99", x"00FE15DC", x"FF5683BF", x"005D5EB7", x"003DD509", x"00C1711B", x"FEEA9A82", x"FFC91DFA", x"FE834DDA", x"FF2B9972", x"FE9A9E16", x"FCEEF4B8", x"FD7251BC", x"FD98D9F8", x"FDDA5B80", x"FEE6291C", x"FEEB91F6", x"FF163BE7", x"000E6CC1", x"FF0C6CB5", x"011696D8", x"004964A1", x"010A0910", x"0086EE55", x"FFF70E6A", x"00CD5BEA", x"FF552595", x"0052816E", x"00804195", x"FF97C859", x"0069D447", x"FEE83A5A", x"FF88753E", x"00C7BC5C", x"00CB73D8", x"FEEE539A", x"00127384", x"FF11788E", x"FF84B942", x"FCD30458", x"FD12DE20", x"FC85BEAC", x"FCB46158", x"FE4C88FA", x"FE67EF6A", x"0145149A", x"0089A82A", x"01C23EB6", x"00FC4B4A", x"01D4D2B8", x"00E77C48", x"01AC8134", x"010EAB60", x"00E088AE", x"FF995A93", x"00B617BA", x"FF0B8DED", x"0084DFAE", x"FFD79516", x"FF206B44", x"FF549CC6", x"FF52B531", x"00C52382", x"FFD4AC6E", x"FF3A1340", x"0003F9C8", x"FD7F5410", x"FD367540", x"FB1A6410", x"FA602CB8", x"F9CC4408", x"FBBC52E0", x"FD7597E8", x"FEBC2C04", x"01538DC4", x"0145CF98", x"01A75AFE", x"032F31A0", x"026176B0", x"002F377E", x"0043B211", x"FFBBA081", x"FF89CCB9", x"FF745D15", x"FF8344B2", x"FF861A89", x"0013CF21", x"01216A88", x"FF8A6F48", x"FFAB742D", x"FF657C9F", x"FFBB83DB", x"FF64B268", x"FD807DD4", x"FD3F8E20", x"FA102890", x"FA2379C0", x"F6DC5020", x"F5E47730", x"F7C14FC0", x"FBF9C7E0", x"FE8F2E4E", x"FE54281E", x"0002E71E", x"0289E650", x"020C3284", x"00EE7F2D", x"001406AA", x"FFEC0002", x"FFBB7D1E", x"FF35FE60", x"FF48983D", x"004BA6C1", x"00B9B79D", x"00E8D618", x"FFC8B530", x"006E2AFF", x"FED5BDF0", x"00252E0E", x"002D6A3B", x"FF7BD21B", x"FD66293C", x"FDD1A67C", x"FA979E10", x"F9CB6540", x"F6E99490", x"F59A4780", x"F8DFB7B8", x"FC21FDDC", x"FEEAD0D0", x"FF171331", x"0070EFF3", x"0094529C", x"01CBCF0E", x"00836C74", x"009F4F2C", x"007A0FDC", x"FEE30FDC", x"FF38D11D", x"00AF76B5", x"010EBB18", x"FEED764C", x"FFC07371", x"FF42A909", x"00BC5616", x"00333ECD", x"000812DD", x"FFB21564", x"FEDB3F80", x"FFC9CDF8", x"FE4C5418", x"FE78FEB6", x"FBE16F58", x"F807C728", x"F8D09C10", x"FD60BF14", x"FFCBAFBE", x"FF80C784", x"FF9AEA8E", x"FFD7B7C8", x"FF1F1216", x"004B9472", x"FE4DA656", x"FF0AA4BF", x"FE770A12", x"FECF63D2", x"FFD7C06E", x"0108685C", x"010E427A", x"004BF0FC", x"0098E883", x"FEFFA970", x"0011E725", x"FFC5754B", x"FE42221C", x"FEE533E0", x"00E305BA", x"01316548", x"00F7AE80", x"00411ABE", x"FE26D0E6", x"FA3E2D98", x"FBF263C0", x"FEDF648E", x"0374B308", x"00858088", x"00835196", x"FF2F15FB", x"FF15EC33", x"FF6EDF21", x"FE8B40D0", x"FEE0704A", x"0076AC20", x"FF016E44", x"008063F3", x"FFB40C9B", x"FF975CF4", x"00A1CF69", x"FFF843B2", x"FE91FA84", x"0081D135", x"FF01378A", x"012A3C82", x"00E9374C", x"03A85D04", x"047E9AE0", x"047335F8", x"027393CC", x"FD01AE14", x"FA733368", x"FE9482B8", x"03787A18", x"03F0A90C", x"02E60088", x"FFF3516B", x"FE1C0B82", x"FDFEA970", x"FF630ECF", x"FE6AF9F2", x"001CB0CF", x"FEA8B736", x"FFFE26A2", x"FF355B8D", x"0067B04A", x"00E7BDCB", x"005960D4", x"FF6C3779", x"FE9AD502", x"FF4B99CF", x"001D9F6F", x"0327B828", x"02F12E2C", x"057E1AA8", x"07B911F8", x"065B5980", x"011761CA", x"FD754EF0", x"FBE8D848", x"0023AA6B", x"04020918", x"04B17470", x"030211E8", x"002FDAD6", x"FF698507", x"FEA44BA0", x"FFBDD30E", x"FF57E5B6", x"FF77AB0E", x"00280039", x"FF118B38", x"00098E98", x"00862CF5", x"FEEBC890", x"FF54F6D0", x"009530D3", x"0006DB98", x"00A88717", x"02AD6D9C", x"03D00FA0", x"067BB4D0", x"06E4CE28", x"07D9D668", x"0740DE58", x"016B806C", x"FE97FB36", x"FE15ED94", x"006F816C", x"057E9588", x"04C21630", x"02CA605C", x"00ADA6F8", x"01AAA64C", x"0080EDC8", x"FED76B3C", x"FFFDF4E3", x"FFB309CA", x"0100D970", x"009E0018", x"FF5247BE", x"0104C5EA", x"FFCAABFE", x"FFB7173A", x"0056A7A7", x"01A57DD4", x"0223AF6C", x"03134ED0", x"05C37DA0", x"080DA890", x"07404CD8", x"0759F6A0", x"0560C450", x"02C7BD38", x"FFF737B6", x"002239FC", x"0313DFC4", x"07744698", x"07CC3A10", x"04D6E140", x"042A2120", x"0304B78C", x"0015AA78", x"00D4D5FC", x"FF21D7F3", x"00AA59DD", x"FF6ADA89", x"0033ABA3", x"FFFC9940", x"0087B6D7", x"002D6913", x"FF2C815C", x"008B25DB", x"0149B38A", x"0194619A", x"03C97BE0", x"05918818", x"06ABFD78", x"06AC8380", x"063E1800", x"055DE6B8", x"0384B340", x"02DF6880", x"02DDD008", x"05083430", x"07DFE3C0", x"06F5E608", x"050A8980", x"03077878", x"0293CF3C", x"002B7E74", x"00B545BC", x"00B0C0DD", x"FECD6F20", x"FF38374B", x"FF13F436", x"004D7654", x"00388659", x"FF68E83C", x"00AE5166", x"006EDE15", x"FF29EF70", x"0180B5C6", x"03231570", x"04FAEB08", x"066F8AC0", x"04D97DF0", x"03243E1C", x"044D9F70", x"02607A94", x"031AB0B4", x"05AB9E80", x"08BCF5F0", x"09626EA0", x"0644C530", x"04C88910", x"019744B2", x"01054BAC", x"FFD1C9C6", x"FFD1D2F0", x"FEB51952", x"FFD23A23", x"00585A7A", x"00D27518", x"FFCD8908", x"010B4B8C", x"FEEB8776", x"FFACCB89", x"002B4E75", x"FFF9A35C", x"00D74DD4", x"00BC8167", x"033BECCC", x"01BE3208", x"014D51D2", x"012D8424", x"00235D59", x"010FBBA4", x"02D3749C", x"06A38F88", x"0713C978", x"05B323E8", x"03613BA4", x"0093852B", x"FEC059BE", x"FE2BD944", x"FD90AD08", x"FF412E3D", x"FE9764E8", x"FF15C5DD", x"FEBE73FA", x"0022233B", x"FFD28D26", x"FF386747", x"00BB87D3", x"00F42CC6", x"FEDC89D2", x"FFE2C028", x"FEF3CFE2", x"FF21992E", x"FFC7F122", x"FEEDF2F4", x"FF4AA0C9", x"FE14CD2A", x"FD29443C", x"FF460791", x"00F4C259", x"03C1C814", x"02E2CE34", x"01AC53EC", x"FF66B370", x"FD6B4FDC", x"FCBC6B50", x"FE7FC2E0", x"FE4864BC", x"FF03268E", x"FE47685C", x"FEF473A4", x"FF629495", x"0002FE61", x"FF2DD9E8", x"002AE434", x"FF43C7E2", x"0029C8B9", x"00C6DC1B", x"FF53F801", x"FF49837F", x"FCBB9324", x"FC85273C", x"FB188330", x"FAE80200", x"FA3897E8", x"FAFB4070", x"FC5E7E84", x"FF3F40A7", x"00BB6335", x"0092F021", x"FF011DE9", x"FF9BB1EE", x"FE8C2CF2", x"FC7F3464", x"FD627E28", x"FE8A90E4", x"FD290958", x"FE12FC4E", x"0033A648", x"FFD56B09", x"005ACCB6", x"FF865178", x"00350BD9", x"00C1CE2A", x"FFB49C46", x"FF633BD7", x"FE1C02B0", x"FE263F76", x"FDD3D4D8", x"FAB149C8", x"FA7DB9A0", x"FAB46F40", x"F997EBB8", x"FAB96A00", x"FC5D18C4", x"FD3D45A4", x"FE6F91DC", x"FDC34FD8", x"FF7581DE", x"FE6F66FE", x"FDF689AC", x"FDAB3320", x"FE9CBC5A", x"FDBF6D80", x"FDDD6FC0", x"FE986D74", x"FEEA3EF6", x"FF5AECEA", x"00E51DEF", x"FF1DA812", x"FF54047A", x"FF1178DC", x"FF68C807", x"FFC99BD3", x"FEC30408", x"FEC05B2A", x"FDE0F900", x"FC0FDCF4", x"FBCFE268", x"FB07CCE8", x"FC107F3C", x"FBED8378", x"FDBF1C28", x"FDD6EFD4", x"FDF51790", x"FF0A4FA4", x"FE34BA1C", x"FEA5C028", x"FFD1A2BE", x"FF8F5FCF", x"002A5673", x"FF3138D7", x"FF4BA466", x"008299BD", x"FFE46777", x"01022F7A", x"FF690AF6", x"FFA001B8", x"000CA3FE", x"009C0A40", x"FEFD3916", x"FF92D546", x"00807558", x"FF660CA8", x"FF251030", x"FD08A450", x"FBFCC040", x"FB900580", x"FBFBFFD0", x"FC57E778", x"FE016DAA", x"FDD3B8AC", x"FD2666B8", x"0032D124", x"00342102", x"01205338", x"00515E01", x"0167982A", x"FF7E0805", x"00FF98DE", x"FF4AC4FA", x"005D9B1D", x"FF88DFFB", x"00B6F7D5", x"FF0A8E17", x"FFC6F46C", x"FFB107BB", x"FF510CEB", x"FF6F9207", x"FFA462FE", x"FFF39D5D", x"00552DF5", x"FEE59FE8", x"FFB67834", x"FDA96074", x"FD732C20", x"FE08150C", x"FE1F09EA", x"FE7BAD12", x"FF201AEF", x"FF1441BD", x"FEF8D888", x"00491738", x"014A36FE", x"00B29CEB", x"01A1E03C", x"01ECF26E", x"01006676", x"0007326E", x"FFE08568", x"FF6EFE9A", x"FFDE2DE0", x"0100C326", x"FF69951D", x"002ECEA7", x"FF295584", x"FFAFDDBE", x"000E6A81", x"FF1008DA", x"001B007C", x"FE9D491A", x"FEE0D584", x"FFEDD800", x"0006B239", x"FEC04C30", x"FE1F0430", x"FD941C08", x"FE0460A6", x"FE329E9C", x"00337649", x"FEF4B126", x"00C90273", x"00BBB604", x"00077A94", x"011153E4", x"00A50F16", x"FFE9D107", x"FF2A8693", x"FFA1AC7B", x"005EE576", x"00FD69EF", x"FF9D44F9", x"FF866989", x"FEE22492", x"00B3C32C", x"011D2662", x"00C472BA", x"FF4410BE", x"00928D43", x"FF1C8FA5", x"FFA9DE0C", x"FF66021A", x"FD67CD88", x"FE02DAD6", x"FDD38B9C", x"FCB50CC8", x"FE8E4F2A", x"FE83C5A2", x"FE9E8308", x"FDD60330", x"FDCB255C", x"FE30BE9A", x"FF9D0E5C", x"FF48D1C2", x"00B58792", x"00E50756", x"000FFBA7", x"FF0FE2F7", x"00740A06", x"0105D21C", x"FFB683D7", x"FF66E1E9", x"FFBB8F49", x"0029DEC5", x"FF249894", x"0095A3E3", x"006151AE", x"FF51B31A", x"FF1E9C74", x"FEC6C8AE", x"00003CDD", x"FF7E1B37", x"FEFB37B4", x"FE80FEEC", x"FEBAF878", x"FFB8351E", x"FF0BDB91", x"FE568094", x"FF998FC3", x"FEF5AFB4", x"FF9CE79B", x"FF18E7F2", x"FFE8E512", x"000DFD9C", x"FF4E82CC", x"00BC0D1D", x"010E3738", x"FF0B4856", x"0054C6DE", x"FF35E3FB", x"FFC5D965", x"008C2580", x"FFFAD8CE", x"00580E78", x"FF9EE936", x"010F1CFA", x"FF6C4857", x"002C5B70", x"000CA5D6", x"00B4C019", x"000647A9", x"0093B5A0", x"001CC110", x"0097C294", x"FFE19539", x"00420BF4", x"0107410E", x"FF9160D1", x"FF82CAAA", x"00D0FBCF", x"006CC537", x"FEEB87A4", x"00680E89", x"FEE10F30", x"FF612804", x"00727EFE"
--  0.020057, 0.016591, 0.020683, 0.009635, -0.013193, 0.014740, -0.016821, -0.021922, 0.033386, 0.029603, -0.025811, 0.029009, 0.007295, 0.008813, 0.034313, -0.001880, -0.011359, 0.022421, -0.009225, -0.008574, -0.014402, 0.035153, 0.017041, -0.005790, -0.000713, 0.002500, -0.021171, 0.010140, -0.027719, -0.001665, -0.006701, -0.014583, 0.033029, 0.009988, 0.016813, -0.024401, 0.004424, 0.008256, 0.016103, -0.013935, -0.011234, -0.031911, 0.019944, 0.021813, 0.014438, 0.016748, 0.020563, 0.033083, 0.011205, 0.012503, 0.010945, -0.020295, 0.008961, 0.010760, -0.028427, -0.010570, -0.022036, -0.022820, 0.024819, 0.028086, -0.005064, 0.010892, -0.008986, 0.004876, -0.010569, -0.025790, -0.027796, 0.017613, -0.015931, -0.040483, -0.015283, -0.053373, -0.015216, 0.015271, -0.004883, 0.003325, -0.036738, -0.009284, 0.019383, -0.026970, -0.017057, 0.024008, 0.010256, 0.016695, -0.033304, 0.022730, -0.007791, 0.007449, 0.028770, -0.033231, 0.008636, -0.036967, 0.016657, -0.006972, -0.023350, -0.051424, -0.031953, -0.068588, -0.043142, -0.018454, -0.069544, -0.046025, -0.018058, -0.009951, -0.007947, 0.025904, -0.012060, 0.008508, 0.018124, -0.007125, 0.023303, 0.023325, 0.015904, -0.008713, 0.031016, -0.020689, 0.011398, 0.007548, 0.023614, -0.033862, -0.006700, -0.046472, -0.025928, -0.043626, -0.095831, -0.079795, -0.075091, -0.067095, -0.034404, -0.033744, -0.028536, 0.001761, -0.029733, 0.034007, 0.008959, 0.032475, 0.016471, -0.001092, 0.025068, -0.020856, 0.010071, 0.015656, -0.012722, 0.012919, -0.034152, -0.014593, 0.024382, 0.024836, -0.033407, 0.002252, -0.029117, -0.015048, -0.099241, -0.091447, -0.108674, -0.102981, -0.053157, -0.049813, 0.039683, 0.016804, 0.054962, 0.030798, 0.057229, 0.028258, 0.052308, 0.033041, 0.027409, -0.012530, 0.022228, -0.029840, 0.016220, -0.004934, -0.027293, -0.020921, -0.021154, 0.024065, -0.005289, -0.024161, 0.000485, -0.078207, -0.087102, -0.153028, -0.175760, -0.193815, -0.133261, -0.079395, -0.039530, 0.041449, 0.039772, 0.051679, 0.099511, 0.074397, 0.005764, 0.008264, -0.008346, -0.014429, -0.017045, -0.015226, -0.014880, 0.002418, 0.035329, -0.014351, -0.010321, -0.018861, -0.008360, -0.018958, -0.078065, -0.085992, -0.185528, -0.183169, -0.285606, -0.315861, -0.257652, -0.125759, -0.045022, -0.052227, 0.000354, 0.079333, 0.063989, 0.029113, 0.002445, -0.002441, -0.008363, -0.024659, -0.022388, 0.009235, 0.022671, 0.028422, -0.006750, 0.013448, -0.036408, 0.004539, 0.005544, -0.016135, -0.081279, -0.068158, -0.168992, -0.193921, -0.283987, -0.324917, -0.222691, -0.120851, -0.033836, -0.028433, 0.013786, 0.018106, 0.056129, 0.016043, 0.019447, 0.014900, -0.034782, -0.024314, 0.021419, 0.033048, -0.033513, -0.007757, -0.023113, 0.022990, 0.006256, 0.000986, -0.009511, -0.035736, -0.006616, -0.053183, -0.047730, -0.128731, -0.249051, -0.224535, -0.081940, -0.006386, -0.015530, -0.012339, -0.004917, -0.027457, 0.009226, -0.053021, -0.029951, -0.047969, -0.037184, -0.004913, 0.032276, 0.032991, 0.009270, 0.018666, -0.031291, 0.002185, -0.007146, -0.054427, -0.034521, 0.027713, 0.037280, 0.030235, 0.007947, -0.057762, -0.179910, -0.126661, -0.035230, 0.107996, 0.016297, 0.016030, -0.025502, -0.028574, -0.017716, -0.045501, -0.035103, 0.014486, -0.031075, 0.015673, -0.009271, -0.012773, 0.019752, -0.000944, -0.044680, 0.015847, -0.031101, 0.036406, 0.028469, 0.114302, 0.140455, 0.139064, 0.076609, -0.093545, -0.173437, -0.044371, 0.108457, 0.123127, 0.090576, -0.001548, -0.059077, -0.062663, -0.019158, -0.049441, 0.003502, -0.041905, -0.000226, -0.024737, 0.012657, 0.028289, 0.010910, -0.018040, -0.043600, -0.022021, 0.003616, 0.098599, 0.091941, 0.171644, 0.241342, 0.198651, 0.034104, -0.079430, -0.127827, 0.004354, 0.125248, 0.146662, 0.094003, 0.005842, -0.018369, -0.042444, -0.008078, -0.020520, -0.016642, 0.004883, -0.029108, 0.001167, 0.016379, -0.033718, -0.020878, 0.018212, 0.000837, 0.020572, 0.083670, 0.119148, 0.202601, 0.215430, 0.245341, 0.226669, 0.044373, -0.043948, -0.059823, 0.013612, 0.171702, 0.148692, 0.087204, 0.021198, 0.052081, 0.015738, -0.036204, -0.000249, -0.009395, 0.031354, 0.019287, -0.021206, 0.031833, -0.006510, -0.008900, 0.010578, 0.051452, 0.066856, 0.096107, 0.180114, 0.251667, 0.226599, 0.229732, 0.168062, 0.086882, -0.001072, 0.004178, 0.096176, 0.232944, 0.243680, 0.151230, 0.130143, 0.094326, 0.002645, 0.025981, -0.027119, 0.020795, -0.018206, 0.006307, -0.000415, 0.016567, 0.005543, -0.025817, 0.016986, 0.040247, 0.049363, 0.118345, 0.174015, 0.208495, 0.208559, 0.195080, 0.167713, 0.109949, 0.089772, 0.089577, 0.157251, 0.246080, 0.217517, 0.157536, 0.094662, 0.080543, 0.005309, 0.022128, 0.021576, -0.037423, -0.024388, -0.028814, 0.009456, 0.006900, -0.018444, 0.021279, 0.013534, -0.026131, 0.046962, 0.098033, 0.155630, 0.201116, 0.151549, 0.098174, 0.134475, 0.074277, 0.097008, 0.177200, 0.273066, 0.293266, 0.195895, 0.149479, 0.049715, 0.031896, -0.005641, -0.005637, -0.040393, -0.005588, 0.010785, 0.025691, -0.006160, 0.032629, -0.033749, -0.010157, 0.005286, -0.000777, 0.026282, 0.023011, 0.101065, 0.054467, 0.040688, 0.036806, 0.004317, 0.033171, 0.088312, 0.207466, 0.221165, 0.178118, 0.105619, 0.018008, -0.039020, -0.057147, -0.076089, -0.023293, -0.044019, -0.028592, -0.039251, 0.004167, -0.005548, -0.024365, 0.022892, 0.029807, -0.035579, -0.003570, -0.032738, -0.027149, -0.006843, -0.033453, -0.022140, -0.059961, -0.088713, -0.022701, 0.029878, 0.117405, 0.090186, 0.052286, -0.018713, -0.080650, -0.102000, -0.046904, -0.053663, -0.030865, -0.053783, -0.032660, -0.019216, 0.000365, -0.025653, 0.005236, -0.022976, 0.005101, 0.024275, -0.021000, -0.022276, -0.102103, -0.108746, -0.153258, -0.159179, -0.180592, -0.156830, -0.113465, -0.023529, 0.022874, 0.017937, -0.031114, -0.012244, -0.045389, -0.109472, -0.081727, -0.045585, -0.088741, -0.060182, 0.006305, -0.005198, 0.011084, -0.014854, 0.006475, 0.023658, -0.009203, -0.019137, -0.059081, -0.057831, -0.067892, -0.165858, -0.172153, -0.165474, -0.200205, -0.164866, -0.113636, -0.086271, -0.048881, -0.069908, -0.016906, -0.048901, -0.063655, -0.072852, -0.043367, -0.070382, -0.066719, -0.043893, -0.033906, -0.020151, 0.027968, -0.027630, -0.020994, -0.029117, -0.018459, -0.006640, -0.038694, -0.039019, -0.066288, -0.123064, -0.130873, -0.155298, -0.122986, -0.127257, -0.070421, -0.067513, -0.063832, -0.029991, -0.056064, -0.042267, -0.005660, -0.013748, 0.005168, -0.025241, -0.022016, 0.015942, -0.003369, 0.031517, -0.018427, -0.011718, 0.001543, 0.019048, -0.031589, -0.013326, 0.015681, -0.018793, -0.026726, -0.092695, -0.125397, -0.138669, -0.125488, -0.114270, -0.062326, -0.067905, -0.089062, 0.006203, 0.006363, 0.035196, 0.009933, 0.043896, -0.015865, 0.031201, -0.022123, 0.011427, -0.014542, 0.022335, -0.029962, -0.006964, -0.009640, -0.021356, -0.017631, -0.011183, -0.001512, 0.010398, -0.034470, -0.008976, -0.073074, -0.079691, -0.061513, -0.058711, -0.047403, -0.027331, -0.028777, -0.032123, 0.008922, 0.040309, 0.021803, 0.051010, 0.060174, 0.031299, 0.000879, -0.003843, -0.017701, -0.004129, 0.031343, -0.018362, 0.005714, -0.026204, -0.009782, 0.001760, -0.029293, 0.003296, -0.043300, -0.035054, -0.002216, 0.000817, -0.039026, -0.058714, -0.075670, -0.061966, -0.056321, 0.006282, -0.032630, 0.024537, 0.022914, 0.000913, 0.033365, 0.020149, -0.002708, -0.026059, -0.011514, 0.011584, 0.030934, -0.012052, -0.014842, -0.034895, 0.021944, 0.034808, 0.023980, -0.022941, 0.017890, -0.027764, -0.010514, -0.018798, -0.081079, -0.062152, -0.067927, -0.102899, -0.045128, -0.046415, -0.043150, -0.067625, -0.068952, -0.056550, -0.012078, -0.022361, 0.022159, 0.027958, 0.001951, -0.029311, 0.014165, 0.031961, -0.008970, -0.018691, -0.008355, 0.005111, -0.026783, 0.018267, 0.011880, -0.021277, -0.027513, -0.038234, 0.000029, -0.015856, -0.031834, -0.046753, -0.039676, -0.008764, -0.029803, -0.051941, -0.012505, -0.032509, -0.012097, -0.028210, -0.002820, 0.001708, -0.021666, 0.022955, 0.032985, -0.029873, 0.010349, -0.024672, -0.007098, 0.017108, -0.000629, 0.010749, -0.011852, 0.033095, -0.018032, 0.005415, 0.001544, 0.022064, 0.000767, 0.018031, 0.003510, 0.018525, -0.003713, 0.008062, 0.032136, -0.013504, -0.015284, 0.025511, 0.013278, -0.033749, 0.012702, -0.035027, -0.019390, 0.013977
--  Sum of weights (converted): FFFFFFFF997B8660
    );

    constant weights_n5 : weight_array := (
     x"009A1E8C", x"FFBDF059", x"00F7A6DE", x"0122C0B8", x"00E423CA", x"FEF3491C", x"FF9594AB", x"0011CCE0", x"00EDCB3C", x"FFCEEC00", x"003D1E32", x"0099FE1C", x"FF66E2F7", x"FF4E83B5", x"01211784", x"FFF9762C", x"00CF051E", x"FEE2B748", x"FF905369", x"00CD4B21", x"FFE3ACC9", x"00628BA0", x"FF0AE834", x"011CC480", x"FF6DF979", x"FFF134D0", x"FF405DE4", x"FF7E319D", x"FF052EA8", x"FEFFEA70", x"FFC43A99", x"FF7EF329", x"00D81E4F", x"FFFE92D8", x"00E35EF2", x"FFCE984A", x"003D3F7D", x"01180CB8", x"FF1CE3F4", x"FF7FF49C", x"00F7D7D9", x"FFBA27E6", x"FFAE4ECF", x"0014C353", x"FF605561", x"0012BD72", x"FF84A7F1", x"005B8043", x"FFC0E154", x"FF9D87E3", x"FF91B673", x"004BFEC9", x"0092D2F3", x"FEF484FC", x"FF33F3B4", x"FEE736CA", x"0088923C", x"00DB6BEE", x"FEE6E52A", x"004BFCA3", x"003B23DC", x"FF62F215", x"003EDC11", x"00E0020E", x"011C0590", x"00788C4E", x"FFB9FF7F", x"FF45BCCE", x"FF72339B", x"FFD56D8F", x"FFAF0F0E", x"009BBC8A", x"FECB4EAE", x"FFF94636", x"FF89667B", x"00003123", x"01008F50", x"FFF59CA9", x"FFC2A23A", x"FF980288", x"FED9EA5E", x"FEF68400", x"007F7A97", x"FF4D5616", x"00A61B45", x"FFAD0D69", x"00698BF2", x"00D55521", x"002BD47D", x"005E8F15", x"00EFC46D", x"FF931A5B", x"00BD3D16", x"FED87BB8", x"00C511B4", x"FF2FEB0F", x"FF72B0DC", x"FFFCE4B6", x"FF674974", x"0061C78B", x"FEF5E51A", x"FF01EE6D", x"00DB4306", x"FF24BAB4", x"00A38E91", x"0106E71E", x"00C429FE", x"FF83CFA9", x"FFF35C3F", x"FEF906C8", x"FF611DAE", x"FFC371A9", x"FF3EB2DF", x"00A8C6DC", x"0099232F", x"FFAAE399", x"FFC82AAE", x"00F1120C", x"FFA42A7F", x"007C08A5", x"003CA276", x"FE974E94", x"FDDA9DF4", x"FFD7B3F2", x"FDBD70F4", x"FEF09DD4", x"FD75D9D8", x"FF0DA332", x"FFEB2D93", x"FFDD6079", x"0150245A", x"FF44C505", x"FFE846D2", x"00CDBE22", x"01FE1C40", x"017B0962", x"0145A624", x"00A62586", x"0111C3D2", x"FFB6CBF0", x"FFA5AE05", x"FFD7D30E", x"00722555", x"FFA178A1", x"003981DC", x"FFCDF3E3", x"FF6ABFBC", x"FFE4DE77", x"FF1478EC", x"FFD98BB6", x"FF3973C7", x"FE8CF61A", x"FFB3D38D", x"FF05F3CF", x"FF9D1701", x"FF767679", x"FFEAD486", x"001E9214", x"0078357F", x"020DDE50", x"037F6A38", x"031BEFBC", x"0344A974", x"03BE1A4C", x"0173E858", x"012D3570", x"FF456426", x"FEF857DA", x"FF555076", x"FFCDE462", x"00613C0D", x"0073C903", x"FED66500", x"FEF442DA", x"FF3D9317", x"FEAB17D8", x"FF4E1EBF", x"00C4E7D9", x"0097E301", x"01BEEFE4", x"018B5E96", x"007A179A", x"FFDDCF79", x"FEE7B4D8", x"FF31E9AC", x"00BA6D11", x"02569FB4", x"036C3CF0", x"037CEB88", x"053198A8", x"04D4EA80", x"05B8D300", x"03C2B63C", x"0271C168", x"01824304", x"0075023F", x"00139A56", x"FF93936A", x"FF08474B", x"FEFCBA1E", x"FE42EED2", x"FFB2342E", x"FE5420E8", x"FF227438", x"FF49F48A", x"00D7CF1E", x"030AA1FC", x"02787640", x"01139A6A", x"00BB7BC2", x"0054EC5E", x"FF461D7D", x"FDE2F9FC", x"FFE998DB", x"000E6C1D", x"015E04B0", x"0416FBD8", x"03897750", x"05271898", x"079F9028", x"07B3E560", x"02A5AE54", x"002192C1", x"FF98658B", x"00E2A2F9", x"00A98067", x"00A889A1", x"0066EAD6", x"FEC4AE28", x"FFA6D9D2", x"FEDA66F0", x"FFC9D2EC", x"00BC9720", x"02303EA4", x"02A5CDC8", x"0247D1B0", x"023C57BC", x"FF756977", x"FF276F7D", x"FF0FABAF", x"FE8E8110", x"FE385508", x"FF1C375D", x"010948E8", x"02684034", x"04042F98", x"060231E0", x"07C48E38", x"06DD9EA0", x"039E6A40", x"020C4690", x"FFEAF558", x"FF8C643D", x"FF273AE0", x"010A4366", x"0041A53E", x"FE83B346", x"FE10845C", x"005B66D0", x"00DEAB20", x"01BA1B50", x"018B44B8", x"0396970C", x"02E7C7FC", x"030FC124", x"0027C521", x"FEDCF020", x"FD5E6E30", x"FE6C9AE4", x"FE795C82", x"FCF76E7C", x"FFC173A4", x"FF9B3295", x"00DF20EC", x"03D6FE80", x"05DA6300", x"06C6CAE8", x"0401E118", x"01D5DD64", x"FF11EFC0", x"00867611", x"FFA074B6", x"FFFF8F0F", x"00876B0A", x"FEB82662", x"00055809", x"FFC8CB04", x"01EB9C4E", x"029641A8", x"043C9370", x"05804518", x"04EB6D28", x"03BC3838", x"04692480", x"00B03E35", x"FF65FEBB", x"FDBD3F0C", x"FB34AA80", x"FBC0D8F8", x"FBF1BA50", x"FC2DA7F8", x"FE0C78C2", x"FF1B598E", x"022E72F4", x"038B2DF0", x"017814BE", x"00A42B8E", x"00A3114F", x"00DF6355", x"005FE9E4", x"006CB9ED", x"FF9648C6", x"FFC54CB0", x"FF19E1D1", x"019AD92A", x"02A59304", x"0280FB30", x"03273FE4", x"0632E4C8", x"05F8A1A0", x"07C14280", x"041C0420", x"0166682C", x"FE3A6274", x"FD29574C", x"F9BC5D30", x"F9C0DDF8", x"F8C5C440", x"FA1A64A8", x"FB28D130", x"FC96AF04", x"FEDE9DF0", x"FF9246BE", x"006F2D9C", x"0096688B", x"01042F18", x"FF9443DA", x"FF16B979", x"FF0FA46D", x"FF5F6AB0", x"00172044", x"000159AE", x"0094EB4E", x"01892552", x"03C09AE8", x"0373F31C", x"079A4728", x"08516F20", x"08436D80", x"059E33C8", x"0103B094", x"FF2FAF4F", x"FBBF64D8", x"FACFDFB0", x"F92FB6D8", x"F9E92058", x"FA513788", x"FA90CC40", x"FB28B138", x"FDA39740", x"FF84972A", x"00C3773F", x"FFD99FEB", x"003223EA", x"FF33B78E", x"FF238527", x"FFC69200", x"0014AEB1", x"FF532D3F", x"FF2B9065", x"00EDB84A", x"02155728", x"0237792C", x"05947498", x"06448158", x"08C26490", x"0771E9A0", x"03701504", x"0174EC2E", x"FCC9B2E0", x"FB7A3560", x"FD23B524", x"FCC74190", x"FCA618CC", x"FCC6D7AC", x"FBFC5FC8", x"FD145EEC", x"FE1480B4", x"FF2DF106", x"001AD22A", x"0047EDAA", x"00068801", x"0023C42D", x"000493EB", x"00C3E318", x"0099213D", x"FFC61FFD", x"FFEB2511", x"FF50BA66", x"0023A590", x"023C50AC", x"030B8A44", x"05D3A2B0", x"0531C5E0", x"033E1E94", x"007AE8BC", x"FE9F35E4", x"FDA04BFC", x"FB722FF0", x"FD0AC254", x"FEDCD73C", x"FE03B5FA", x"FF333430", x"FE0F453C", x"FC921610", x"FDEA1124", x"FDF0394C", x"00D5BDCE", x"00847B57", x"006FED14", x"00E10F52", x"00DF38E1", x"011FD292", x"00700D47", x"FEE49E70", x"FFC14990", x"FE3DDB5A", x"FD35B6B0", x"FE319214", x"01596F00", x"01A05A90", x"01FFDE30", x"006DCAB4", x"FF7E313C", x"FBE87310", x"FC2816D4", x"FC7A1A6C", x"FD36FF18", x"00153401", x"FFF195AA", x"FF905926", x"FFA1E67B", x"FE7D6B26", x"FEB3F418", x"FE711564", x"FFDAC8F0", x"FF6F8DEE", x"00A86CF4", x"00FE6DE6", x"FEEEBD44", x"FF51EA1C", x"01129D8E", x"FF2B2519", x"FF91CD05", x"FEC2D94A", x"FC3A581C", x"FAEB8C78", x"FCABD3F4", x"FCFC8CBC", x"FD93461C", x"FD0FE444", x"FD488048", x"FB902220", x"FCD803B8", x"FD69B2A4", x"FEF4CCB6", x"FEFFF9F2", x"002D179E", x"FF940EAD", x"FEC17FA4", x"FFDF9C9C", x"FFA9AEC9", x"00349DFD", x"FFD54CF0", x"FFEECB18", x"FFF3293A", x"009E093E", x"FF353DDD", x"0037B896", x"00925A15", x"0069DFB7", x"FEFB787E", x"00914609", x"FD1DE1E4", x"FC4BEFB8", x"FB6EEAA8", x"FA0FAB70", x"FAEDE368", x"FA202778", x"FBA540A0", x"FCA35CC8", x"FCE431D4", x"FEBC6330", x"006AABC6", x"0053F2B3", x"01CB234A", x"FFCA72AE", x"00C1857C", x"00CC08EA", x"012522C2", x"FFAA061D", x"FED6492C", x"FF8DD57D", x"00D84BF2", x"00197E6F", x"01175868", x"FF208420", x"FF28C8EA", x"00764139", x"00D00838", x"0180B816", x"01F84A0E", x"FDC07F10", x"FB337FA0", x"FB4D5020", x"FAB6A688", x"FBF200F0", x"FD2F2B3C", x"FF2E106E", x"FFF47758", x"00A246D8", x"FFDEF32D", x"0069CD86", x"01EAAD56", x"00720AFA", x"002BC84A", x"002E4D9F", x"FF6FA646", x"FF78AFF2", x"00ECAB35", x"00326D0B", x"0035DBD7", x"0073FBD8", x"00B138C6", x"00BE59E4", x"00983281", x"003E8C03", x"01B163CA", x"043FF1D8", x"035C6DD4", x"0230B0F8", x"FF4B610A", x"FDB01160", x"FFBA21A1", x"FE956B14", x"FF4C8E46", x"FEEDF69C", x"FEE37C00", x"FFFFD141", x"0111F3A8", x"0028E0EA", x"0112F2D6", x"003DEA41", x"010D2140", x"01762A90", x"00465945", x"FFD0124D", x"00B008F2", x"FF3FDF73", x"FFC3D7D1", x"FF0C6898", x"00CC575E", x"0055B291", x"FF453FF8", x"0054848E", x"018160B0", x"038E8F10", x"03B51A08", x"047C3778", x"04935668", x"033860AC", x"015F091E", x"01BE2D70", x"FFB58B63", x"FFBE6B9F", x"FFFF9C78", x"0015D104", x"004D0E67", x"01F211D6", x"02063F00", x"01F54936", x"00485859", x"00FDC356", x"00AE367D", x"FFF4310F", x"FFBD60B3", x"FF948E33", x"0064D469", x"008B0764", x"FFC6C000", x"00D9680F", x"FFC4F046", x"FFDF9DE5", x"FFF9B18C", x"0106AE84", x"036D1E30", x"0490B810", x"05204588", x"035F7384", x"0279378C", x"00652EB3", x"FFD10B5F", x"FFF2C4F8", x"00D8C57A", x"FFEE7761", x"019B86D0", x"02A05418", x"01031650", x"02469E4C", x"017C3ACE", x"FFF27D2F", x"00A1FF47", x"FF5CBD63", x"003D2F31", x"FEF9A3B6", x"0112EA52", x"FF832B1B", x"00BB17A9", x"FF3E8ABB", x"FEE1491A", x"00367B07", x"002A1F94", x"FFDAD0CA", x"004EE144", x"025E3CF4", x"02C3DAE8", x"03D23704", x"034045BC", x"03212000", x"02FF758C", x"0115DE18", x"02D3A590", x"036B2788", x"02A1F0C8", x"0125164A", x"0104AEE0", x"01B9FE20", x"019CB6D2", x"0108E69E", x"004E6289", x"FF5B7CD5", x"FF07F72F", x"FF5B10B6", x"00022CBB", x"00269069", x"00E012C1", x"FF2A21A9", x"0089D661", x"00E00958", x"FEC84C3C", x"FF2D114E", x"FFF4489D", x"01673BBA", x"0306E1E8", x"02DDDD8C", x"03D22168", x"0400BEC0", x"03B5C93C", x"01C526D6", x"01CBBCA2", x"0226B060", x"0174F214", x"00F6E231", x"01953DD0", x"0169B04A", x"FFBCE3E4", x"FF828785", x"002B4680", x"0032044E", x"00BB735B", x"00693FA4", x"005B2B2B", x"00600C82", x"00D9D3F5", x"00AD95D9", x"FFE0AFE3", x"FF1F07B6", x"009D2B97", x"FFC49979", x"FF474465", x"0027194A", x"01DD4534", x"00E1F035", x"01D1CBD8", x"02B0CD50", x"03183AD0", x"01C1AB72", x"00589CDC", x"FFE185FF", x"FFC7FBD0", x"002C59CA", x"FF26647F", x"00E52D79", x"00388848", x"FF34DB61", x"00AADFC1", x"001858D8", x"011CC924", x"FFFA135A", x"FFFC2447", x"FEE5A1FC", x"FF0E56BF", x"0001023B", x"00FAD711", x"FF4978FA", x"0021D9EA", x"FF0EEE1B", x"FEF9C460", x"FF7341C8", x"FF485C4C", x"FF328FCB", x"FFF84383", x"00309DDB", x"00CE5C03", x"0063C13E", x"FFBFE892", x"FF73E590", x"FF8535EE", x"FECD2D10", x"00904DF9", x"00D82700", x"FEEE89DA", x"FEFA0EAA", x"FEFEF0DE", x"FFDB7F81", x"FFFF39CB", x"FF40F3F2", x"00A1AB13", x"0013447D", x"FF6BE8A2", x"FEE4F740", x"00E3C260", x"011F10C0", x"0013921C", x"FF6419C0", x"009BDA47", x"007D0C8C", x"FF9F40F7", x"00D51D3B", x"FEEAC4D0", x"FF9E839D", x"00A19290", x"FEE80B32", x"FF5F6D55", x"FF3ED2F2", x"FF49C6AC", x"00C79CB7", x"009111BF", x"FEE94AB8", x"FF4BBD23", x"FFFD91EF", x"FFA06CE3", x"FF5EC7E3", x"FEE06198", x"00D7C75A", x"00A3CE90", x"0054E42B", x"FFBE2870", x"FEE46784", x"FFEDAEFC", x"006FD712", x"FFAAC169", x"00E58278", x"00415E7C", x"FFEEFC07", x"00707174", x"009627A6", x"FF28DE8A", x"0053A3CA", x"FEE91A38", x"FFB09EA6", x"FF92EBDD", x"00D1709D", x"FED8A634", x"005D2299", x"FEEF47E0", x"007C2F8A", x"004680A3", x"FF8BF676", x"005651E8", x"0118CD36", x"00B21EA3", x"FEF509BC", x"FFB42D8E"
--  0.018813, -0.008064, 0.030231, 0.035492, 0.027849, -0.032802, -0.012991, 0.002173, 0.029028, -0.005991, 0.007461, 0.018798, -0.018691, -0.021666, 0.035290, -0.000798, 0.025271, -0.034825, -0.013632, 0.025060, -0.003458, 0.012029, -0.029919, 0.034762, -0.017825, -0.001806, -0.023393, -0.015845, -0.030617, -0.031260, -0.007296, -0.015753, 0.026382, -0.000174, 0.027755, -0.006031, 0.007477, 0.034186, -0.027723, -0.015630, 0.030254, -0.008526, -0.009972, 0.002535, -0.019491, 0.002288, -0.015057, 0.011170, -0.007705, -0.012020, -0.013463, 0.009277, 0.017923, -0.032651, -0.024908, -0.034276, 0.016671, 0.026785, -0.034315, 0.009276, 0.007219, -0.019172, 0.007673, 0.027345, 0.034671, 0.014715, -0.008545, -0.022737, -0.017309, -0.005197, -0.009881, 0.019011, -0.037682, -0.000821, -0.014478, 0.000023, 0.031318, -0.001268, -0.007491, -0.012694, -0.035899, -0.032408, 0.015561, -0.021810, 0.020277, -0.010125, 0.012884, 0.026042, 0.005350, 0.011543, 0.029268, -0.013293, 0.023100, -0.036074, 0.024056, -0.025401, -0.017250, -0.000379, -0.018642, 0.011936, -0.032484, -0.031014, 0.026765, -0.026766, 0.019965, 0.032093, 0.023946, -0.015160, -0.001543, -0.032101, -0.019395, -0.007392, -0.023596, 0.020603, 0.018694, -0.010390, -0.006816, 0.029428, -0.011210, 0.015141, 0.007402, -0.044030, -0.067063, -0.004919, -0.070625, -0.033128, -0.079364, -0.029585, -0.002542, -0.004226, 0.041033, -0.022855, -0.002896, 0.025115, 0.062269, 0.046269, 0.039752, 0.020282, 0.033419, -0.008936, -0.011025, -0.004904, 0.013934, -0.011539, 0.007020, -0.006109, -0.018219, -0.003312, -0.028751, -0.004694, -0.024237, -0.045293, -0.009299, -0.030523, -0.012074, -0.016789, -0.002584, 0.003732, 0.014674, 0.064193, 0.109304, 0.097160, 0.102132, 0.116956, 0.045399, 0.036769, -0.022779, -0.032185, -0.020836, -0.006117, 0.011869, 0.014134, -0.036329, -0.032683, -0.023734, -0.041615, -0.021714, 0.024036, 0.018541, 0.054558, 0.048263, 0.014904, -0.004174, -0.034216, -0.025157, 0.022757, 0.073074, 0.106963, 0.108999, 0.162304, 0.150991, 0.178812, 0.117519, 0.076386, 0.047151, 0.014283, 0.002393, -0.013235, -0.030239, -0.031650, -0.054329, -0.009497, -0.052230, -0.027044, -0.022222, 0.026344, 0.095048, 0.077205, 0.033643, 0.022886, 0.010367, -0.022691, -0.066043, -0.002735, 0.001761, 0.042727, 0.127806, 0.110531, 0.161022, 0.238228, 0.240710, 0.082725, 0.004098, -0.012647, 0.027666, 0.020691, 0.020573, 0.012563, -0.038491, -0.010882, -0.035840, -0.006613, 0.023021, 0.068389, 0.082740, 0.071267, 0.069866, -0.016917, -0.026436, -0.029337, -0.045104, -0.055624, -0.027806, 0.032383, 0.075226, 0.125511, 0.187768, 0.242744, 0.214553, 0.113088, 0.063998, -0.002569, -0.014112, -0.026461, 0.032503, 0.008013, -0.046423, -0.060484, 0.011157, 0.027181, 0.053968, 0.048251, 0.112133, 0.090794, 0.095673, 0.004855, -0.035530, -0.082223, -0.049243, -0.047685, -0.094796, -0.007635, -0.012305, 0.027237, 0.119994, 0.182909, 0.211767, 0.125229, 0.057357, -0.029060, 0.016414, -0.011663, -0.000054, 0.016531, -0.040021, 0.000652, -0.006739, 0.060011, 0.080842, 0.132395, 0.171908, 0.153739, 0.116726, 0.137835, 0.021514, -0.018799, -0.070649, -0.149821, -0.132709, -0.126742, -0.119427, -0.060978, -0.027911, 0.068170, 0.110740, 0.045908, 0.020040, 0.019906, 0.027269, 0.011708, 0.013272, -0.012905, -0.007166, -0.028091, 0.050152, 0.082712, 0.078245, 0.098541, 0.193713, 0.186601, 0.242341, 0.128420, 0.043751, -0.055373, -0.088703, -0.195756, -0.195207, -0.225859, -0.184278, -0.151267, -0.106606, -0.035325, -0.013394, 0.013572, 0.018360, 0.031761, -0.013151, -0.028476, -0.029341, -0.019602, 0.002823, 0.000165, 0.018179, 0.047991, 0.117261, 0.107904, 0.237583, 0.259941, 0.258231, 0.175562, 0.031700, -0.025429, -0.132886, -0.162125, -0.212926, -0.190292, -0.177586, -0.169824, -0.151283, -0.073780, -0.015065, 0.023861, -0.004684, 0.006121, -0.024937, -0.026914, -0.007010, 0.002525, -0.021097, -0.025932, 0.029019, 0.065105, 0.069272, 0.174372, 0.195862, 0.273730, 0.232655, 0.107432, 0.045523, -0.100379, -0.141332, -0.089391, -0.100677, -0.104725, -0.100727, -0.125443, -0.091263, -0.059997, -0.025642, 0.003274, 0.008780, 0.000797, 0.004366, 0.000559, 0.023912, 0.018693, -0.007065, -0.002546, -0.021395, 0.004351, 0.069863, 0.095159, 0.182084, 0.162326, 0.101333, 0.015004, -0.043065, -0.074183, -0.142311, -0.092437, -0.035542, -0.062047, -0.025000, -0.060636, -0.107167, -0.065177, -0.064426, 0.026091, 0.016172, 0.013663, 0.027473, 0.027249, 0.035135, 0.013678, -0.034592, -0.007655, -0.054949, -0.087193, -0.056449, 0.042167, 0.050824, 0.062484, 0.013402, -0.015846, -0.127875, -0.120106, -0.110095, -0.087037, 0.002588, -0.001760, -0.013629, -0.011487, -0.047190, -0.040533, -0.048696, -0.004543, -0.017633, 0.020560, 0.031058, -0.033357, -0.021251, 0.033522, -0.025983, -0.013452, -0.038715, -0.117878, -0.158746, -0.104025, -0.094171, -0.075772, -0.091810, -0.084900, -0.138656, -0.098631, -0.080847, -0.032617, -0.031253, 0.005504, -0.013177, -0.038880, -0.003954, -0.010537, 0.006423, -0.005212, -0.002100, -0.001567, 0.019292, -0.024751, 0.006802, 0.017865, 0.012924, -0.031803, 0.017734, -0.090102, -0.115730, -0.142710, -0.185587, -0.158461, -0.183575, -0.136078, -0.105058, -0.097144, -0.039503, 0.013021, 0.010248, 0.056047, -0.006537, 0.023623, 0.024907, 0.035783, -0.010495, -0.036342, -0.013936, 0.026403, 0.003112, 0.034100, -0.027281, -0.026271, 0.014435, 0.025395, 0.046963, 0.061559, -0.070252, -0.149964, -0.146812, -0.165204, -0.126709, -0.087992, -0.025627, -0.001408, 0.019809, -0.004034, 0.012915, 0.059897, 0.013921, 0.005345, 0.005652, -0.017621, -0.016518, 0.028890, 0.006156, 0.006575, 0.014158, 0.021634, 0.023236, 0.018579, 0.007635, 0.052904, 0.132806, 0.105033, 0.068444, -0.022048, -0.072257, -0.008529, -0.044260, -0.021905, -0.033452, -0.034731, -0.000022, 0.033441, 0.004990, 0.033563, 0.007558, 0.032853, 0.045675, 0.008587, -0.005851, 0.021489, -0.023453, -0.007343, -0.029735, 0.024944, 0.010461, -0.022797, 0.010317, 0.047043, 0.111152, 0.115857, 0.140163, 0.142986, 0.100632, 0.042851, 0.054465, -0.009089, -0.008005, -0.000047, 0.002663, 0.009406, 0.060800, 0.063262, 0.061192, 0.008831, 0.030977, 0.021266, -0.001441, -0.008133, -0.013116, 0.012308, 0.016971, -0.006989, 0.026539, -0.007210, -0.003953, -0.000770, 0.032066, 0.107070, 0.142666, 0.160189, 0.105402, 0.077297, 0.012351, -0.005732, -0.001615, 0.026461, -0.002140, 0.050235, 0.082071, 0.031627, 0.071120, 0.046415, -0.001649, 0.019775, -0.019929, 0.007469, -0.032026, 0.033559, -0.015238, 0.022838, -0.023615, -0.034999, 0.006650, 0.005142, -0.004539, 0.009629, 0.074004, 0.086408, 0.119411, 0.101596, 0.097794, 0.093684, 0.033919, 0.088336, 0.106830, 0.082268, 0.035777, 0.031822, 0.053954, 0.050380, 0.032337, 0.009568, -0.020082, -0.030278, -0.020134, 0.000265, 0.004708, 0.027353, -0.026107, 0.016826, 0.027348, -0.038050, -0.025749, -0.001430, 0.043852, 0.094590, 0.089583, 0.119401, 0.125091, 0.115941, 0.055316, 0.056120, 0.067223, 0.045526, 0.030137, 0.049468, 0.044151, -0.008192, -0.015316, 0.005283, 0.006106, 0.022882, 0.012848, 0.011129, 0.011725, 0.026590, 0.021190, -0.003822, -0.027462, 0.019186, -0.007251, -0.022550, 0.004773, 0.058261, 0.027580, 0.056860, 0.084082, 0.096708, 0.054891, 0.010817, -0.003720, -0.006838, 0.005414, -0.026563, 0.027976, 0.006901, -0.024798, 0.020859, 0.002972, 0.034764, -0.000723, -0.000471, -0.034469, -0.029500, 0.000123, 0.030620, -0.022281, 0.004132, -0.029427, -0.032011, -0.017181, -0.022417, -0.025078, -0.000944, 0.005935, 0.025190, 0.012177, -0.007824, -0.017102, -0.014989, -0.037454, 0.017615, 0.026386, -0.033382, -0.031975, -0.031379, -0.004456, -0.000095, -0.023321, 0.019735, 0.002352, -0.018078, -0.034550, 0.027803, 0.035042, 0.002389, -0.019031, 0.019025, 0.015265, -0.011810, 0.026015, -0.033842, -0.011900, 0.019723, -0.034174, -0.019601, -0.023581, -0.022244, 0.024367, 0.017709, -0.034022, -0.022005, -0.000297, -0.011667, -0.019680, -0.035110, 0.026340, 0.019996, 0.010363, -0.008037, -0.034619, -0.002236, 0.013652, -0.010406, 0.028016, 0.007980, -0.002077, 0.013726, 0.018329, -0.026261, 0.010210, -0.034045, -0.009690, -0.013315, 0.025566, -0.036054, 0.011369, -0.033291, 0.015159, 0.008606, -0.014165, 0.010537, 0.034278, 0.021743, -0.032588, -0.009256
--  Sum of weights (converted): 000000009FD127B4
    );

    constant weights_n6 : weight_array := (
     x"01096320", x"002D43AB", x"002411CD", x"0014DFCD", x"FF9922DB", x"FFB37749", x"00136AB2", x"00DC3BE3", x"FFAD8A0B", x"FFB36FA2", x"0037B19E", x"FF94EAD0", x"01007DA8", x"00DE78C7", x"000BCA99", x"FF42C82A", x"0051E18B", x"00F81D95", x"00606282", x"007AA225", x"FF65234B", x"FEDFC92C", x"FF91FC2B", x"00095999", x"0103F0EE", x"003D1660", x"FFCA5DA3", x"FFB67BE7", x"FFC80F25", x"FF62AD02", x"FF8583C2", x"00365A84", x"00C636D9", x"00F8C8E5", x"0076549A", x"FF44B1C0", x"0123F206", x"013724D6", x"FFD26E6D", x"00425CE7", x"014C4380", x"FFCBBDCB", x"00AB187E", x"004ECCF3", x"00BF4EFC", x"0085571A", x"013BE842", x"010AA406", x"FF4745CE", x"00B8BA88", x"FFCA8E18", x"FF686211", x"0031124D", x"FFD82D67", x"FF4156E6", x"FEFDC0D2", x"FF5CF259", x"001E1F3D", x"00B2507C", x"00AC61F3", x"005187D3", x"0116C828", x"FF125D1D", x"FF7559D2", x"00D0A7DC", x"FF83EAB1", x"020CDFC0", x"016EF97A", x"013220B8", x"02DCB428", x"028486F4", x"02DC936C", x"02BBDBA4", x"01A3C7A8", x"02BBAFEC", x"01927704", x"0114087C", x"010BCBC2", x"FF7F1890", x"FF77D335", x"011E50CA", x"FF40B9CA", x"009E1643", x"00B0D237", x"FF1279CF", x"FFDE7817", x"FFFCD78B", x"00D9C072", x"FFB30259", x"010BF06E", x"FF2563BE", x"00BBE9D9", x"011C1870", x"0069ADAA", x"00F48AB8", x"00FA0562", x"025413F4", x"02F77BE4", x"02EABED0", x"04D9C000", x"045187E0", x"04D4EC38", x"05CC29F0", x"04B54FD8", x"03FD958C", x"02F7C2F0", x"008BB2E9", x"00A22C49", x"014D2946", x"FF540C10", x"0028CB73", x"00D9547C", x"00204DC7", x"FFBE6572", x"00699DE9", x"FF0D9C5A", x"00F0D08F", x"00DE36B7", x"FFA90BB6", x"FF9E4027", x"000A4819", x"019D20F0", x"004531D6", x"00C7CC4C", x"FF618DF9", x"0128F964", x"01F6777E", x"026553D4", x"0345C554", x"04AE84B0", x"060D86E8", x"05471940", x"037847E0", x"01B21894", x"025D5AA4", x"00540FD7", x"00FC16B7", x"FFD2C7EE", x"0003FDF9", x"FF1ABC98", x"FF908A87", x"001823CB", x"FEE56C4A", x"FFBE902F", x"00A0D9C2", x"009D6971", x"0085E4E6", x"FF440E08", x"FFF4DF0E", x"FEF42E90", x"004F7AA5", x"FF319566", x"FFE3341F", x"FE8023AC", x"0001561A", x"0019D748", x"0193942A", x"019CB21E", x"015D32A4", x"013F0C2E", x"00531EFF", x"00F93628", x"FF6F5CC3", x"FFBD7C99", x"009A739F", x"0105A0B6", x"FFB5C4B3", x"00CCA09D", x"FFE9D47C", x"FFC5735F", x"FFDCC2A1", x"FF6C470D", x"002BA73E", x"FFA55E01", x"FED57C30", x"001F6820", x"FEE0FC86", x"FE8655BC", x"FF27E780", x"FE474E18", x"FD8725DC", x"FC93E85C", x"FD07716C", x"FD0E6D78", x"FEDF90E6", x"FE125AAE", x"FEA0CF40", x"FE92AD04", x"FE1F39D0", x"FE18A1F0", x"FE1774E2", x"FF4A1B3C", x"FE7054BA", x"FF353F3C", x"00DA5072", x"FFC819A1", x"00EC062C", x"00AD2C72", x"FFC0C57C", x"FEFBB216", x"00ADFC9E", x"FF8E256C", x"003324A4", x"FE2D8E28", x"FF58D72B", x"FE004EF8", x"FE32E7C8", x"FCFDC378", x"FC6DA884", x"FCE0D704", x"FE2882B0", x"FD644AD8", x"FC26EA08", x"FC35A734", x"FA781908", x"F9EB73A0", x"FC123AC0", x"FD1E0DF0", x"FE3F715C", x"FF06E1FB", x"00148E90", x"FF1D3AC8", x"00103B40", x"FF951F5E", x"FFD908E6", x"00E715E4", x"FF13D0D3", x"007F483E", x"FF01C30A", x"FF41D9A7", x"FECC9EF2", x"FE95941E", x"FF3A8B39", x"FE606912", x"FF3AEEE7", x"FD9F63FC", x"FE3128F8", x"FD34CC98", x"FCE8EC1C", x"FD9DD1C8", x"FA610350", x"F85EC360", x"F80B0AF8", x"F8AB5FD8", x"FA603D40", x"FB0F4D40", x"FC3DB994", x"FE5CBDB6", x"FF342786", x"00688D73", x"FFFC8EAB", x"FFB17E39", x"FFC16103", x"FFC3AAA0", x"FF9BCC32", x"FF7078F8", x"FF440D9E", x"FF84D983", x"FF80A993", x"003BF1D1", x"FE7F69B2", x"FFE779BF", x"FE871D6A", x"FD66547C", x"FF6AF644", x"FE88FE3A", x"FE56FB02", x"FC93A3A0", x"F9A37A00", x"F8760C28", x"F6CEA8C0", x"F94571D8", x"FAC74A40", x"FC55FB1C", x"FC7A2B14", x"FE45CBD6", x"FF2CA94D", x"007CCFEA", x"FF28B73E", x"FEF05B74", x"FEF6F9DC", x"00258762", x"FF17E09F", x"FF9DE3F7", x"FF077F0C", x"FF7AA3F8", x"FE925A06", x"009B537F", x"FEFE8862", x"FEF78F64", x"FFBF87F0", x"FE686CE4", x"007D153A", x"00633CCC", x"FE07AAF2", x"FBFB1938", x"F8B30AB0", x"F8F04178", x"F8CE8088", x"FAB63298", x"FCB8F5EC", x"FE585D00", x"FDB8953C", x"FE0B7210", x"FE9A3162", x"FFE715D3", x"0055F309", x"0095CA75", x"007EE4A7", x"011ACBCA", x"FF1B9FDA", x"FEF1867C", x"FF3DF835", x"006A2B67", x"FEF3F96A", x"01494690", x"00BD1811", x"0127F850", x"0158BDCA", x"01C58252", x"02EE9F50", x"00D497DD", x"FCF9322C", x"FB03F960", x"FB984250", x"FB3CFB08", x"FBA6A508", x"FCA6DF10", x"FDD6A544", x"0076ABF2", x"FFA987CE", x"01E0A918", x"00266CD4", x"FF253142", x"FF7F3F83", x"FF4AE687", x"FF01BF89", x"001C5501", x"FFB8FD1B", x"FF59F2F3", x"FF62C704", x"FF7A70AA", x"00BE1F2B", x"FFE99EF3", x"00FD53C5", x"00EB3C62", x"00123807", x"0337F73C", x"02052BFC", x"00F2A2AB", x"FD6B2884", x"FC109724", x"FE40B020", x"FD162898", x"FE1DFCD0", x"FE05A818", x"FFC5F8FA", x"02552724", x"03703614", x"01ACDC64", x"00A82FF9", x"FF622F2F", x"FFD0DBEA", x"FF0B82DE", x"FF186C3A", x"FFBF5328", x"0116BC9E", x"0016656A", x"FF198A99", x"008376F8", x"015528C4", x"01CCF998", x"0170DFC4", x"01783112", x"03105AFC", x"03BD63D4", x"02D577B4", x"FFB12987", x"FD52D86C", x"000AC943", x"0066EB16", x"010779F2", x"009C9DE4", x"012B6490", x"0242A694", x"03EB1E38", x"031A4E04", x"02DD6AE8", x"01809794", x"FF88AA9D", x"00BD039D", x"0016D36F", x"FFB5D58E", x"FF7CA9D9", x"FEFA808E", x"FFFE44CE", x"007D1088", x"006764A1", x"016772CA", x"021933C4", x"02493BB8", x"0286B008", x"029E59B4", x"047B4420", x"00750291", x"FE227F14", x"0025F682", x"023FBF18", x"018FB93A", x"01437D6A", x"FE95B708", x"00B29F00", x"027EE8D0", x"03A976B4", x"035A4B08", x"028E0E78", x"02A796AC", x"006F76DD", x"FF5DD208", x"01191A80", x"FFC2E80A", x"FFC9DB91", x"004A2017", x"00D01169", x"FED640DE", x"FF687F4D", x"FFE44DAB", x"00EEA0D6", x"02101D50", x"03853098", x"05385288", x"031EEBF4", x"01CDE6EC", x"00F52484", x"0189F790", x"0237E898", x"01A3C42A", x"FEEE92A6", x"00688B86", x"0057771D", x"024631E0", x"042AEB10", x"041716F8", x"022807C0", x"0079D7CD", x"FF03BE91", x"FED936A0", x"FFBEBCEE", x"FF1CD9E1", x"FFE26458", x"FF620C34", x"0074C97A", x"FFFD0DEC", x"0009A357", x"FF348789", x"00B225B8", x"032F75A8", x"045124D0", x"069CE9D8", x"03C31D8C", x"02B676B4", x"0041DE41", x"009699DD", x"00786836", x"FE9111CA", x"FDFE59A8", x"00B1F9B2", x"02477220", x"032BFFE0", x"03248980", x"02ACCFE0", x"011C0A2C", x"01BBC582", x"FF39B1D1", x"FECC9306", x"00F24B42", x"FFE86790", x"00C477C2", x"FF99A714", x"00A263F2", x"FE30F7B6", x"FF43E32B", x"000E1BF8", x"0133C7E2", x"04082C88", x"0565CFD8", x"060F5BE8", x"06901898", x"022FBC70", x"0182CEA2", x"FF740C47", x"FE501562", x"FDEF7A6C", x"FF408C4B", x"00B5CD81", x"02722FB8", x"020F3C84", x"01DC083A", x"00DA45D9", x"0020E07A", x"FF994E77", x"00ADA02A", x"FF08DFB9", x"FF1D9F9B", x"FF11CD23", x"01119D78", x"FFD512FE", x"FF5EC1DC", x"FF7FC003", x"FD6CDE40", x"FE129AC8", x"0166AA42", x"0394F564", x"04CFAA88", x"07A337A8", x"0789F740", x"0557A7F8", x"0194590C", x"011AD228", x"FFDF0660", x"FFDEF350", x"02F160B0", x"02E7A7F0", x"03C9926C", x"01E1433E", x"01E2CA68", x"009E230E", x"FEDDEEAC", x"FF0D4422", x"FFAEC090", x"FF425DFC", x"00241AC0", x"009A7EE4", x"00220096", x"FED8EBDA", x"FFA70A08", x"FE56248A", x"FE3E320A", x"FCEEBE88", x"FE4F1372", x"01521BEE", x"05082678", x"074998C8", x"086E4C90", x"06AC2190", x"0309FA50", x"026F06C8", x"02F3210C", x"044C2450", x"053BE3C8", x"04ACC4F0", x"03D95260", x"01E925E2", x"0058ED61", x"00AC64C5", x"001A8727", x"FFE9C013", x"00771922", x"0075298A", x"00FF4F39", x"00FE81EA", x"FF1152FF", x"FEE46A90", x"FF1BFF64", x"FFD7DF54", x"FF0359E3", x"FD6B0734", x"FCFE04B8", x"FE9F7E12", x"0248B4BC", x"0646C948", x"07BE9298", x"07376D98", x"080C2B40", x"075E2390", x"059A8080", x"0501ACA8", x"050EDFA0", x"024DE6B4", x"026A2644", x"FFFD4FED", x"FF2B5BE2", x"FE3C5D3C", x"FDF6C25C", x"FFB37059", x"FF64A39A", x"FF4BA7A4", x"00E9354C", x"00364047", x"FFB17D4B", x"FEECC450", x"FF2C3525", x"FEE9A6A8", x"FEDA71D6", x"FC5D3EEC", x"FDB5B3E0", x"FE727D02", x"FEF7D60C", x"FFEA031F", x"03E71F48", x"05608A78", x"06DECEC8", x"05EE4708", x"0528D9D8", x"02D34D10", x"01AF52FE", x"00A2F754", x"FE401FAC", x"FEC5B88C", x"FF965ABC", x"FFC71E94", x"FF75A865", x"FF7D94E6", x"005EA890", x"FEFBB5DC", x"FFA7E118", x"00FDC3FC", x"0025A647", x"FFF9ABE6", x"FF036190", x"FEE7A74A", x"FF381FE0", x"FD49DB00", x"FCE529AC", x"FBE43DC8", x"FC5B34E4", x"FC8C3ECC", x"FBF1FD90", x"FE7D11AC", x"FE880472", x"FDE4FF1C", x"FEFB1954", x"FCF51FDC", x"FC722BC0", x"FDA1BE40", x"FD46D1F8", x"FDF2C1AC", x"FDE93A08", x"FEFD9412", x"00817D46", x"FECD4B02", x"FF2E96EA", x"FFBF086A", x"FF1873CD", x"0036C3F2", x"FFC5DC50", x"00DCABE1", x"FED56FF0", x"FFE9900D", x"00238D64", x"FF53B907", x"FE19BADE", x"FE7BF8C2", x"FB7969F8", x"FC47BF14", x"FAB2EFA0", x"FA950EA0", x"FAFD4470", x"FAA0FDD0", x"FB4927E8", x"FBB8BD20", x"FBBEBB98", x"FE3D7110", x"FF57C2FF", x"FF71BFA2", x"FF2A9D1C", x"FE9D5558", x"FFC99539", x"00373164", x"FF160CA1", x"00F845BF", x"FFF84BAC", x"004FE892", x"01021A26", x"007EF608", x"FF6082A8", x"00640C00", x"008FD70C", x"004B4037", x"FEE43E78", x"FF17BD10", x"FD9EF654", x"FDBB73E4", x"FC898D48", x"FDB623FC", x"FE169514", x"FC0919B8", x"FCFF8C5C", x"FD83D8AC", x"FDA21F04", x"FFE297AF", x"FE4E371C", x"FEDFAEC6", x"FEBBC0FE", x"FFD30563", x"FF127384", x"FF348C28", x"01221B02", x"0082ABB0", x"007C1F29", x"00CF7D9A", x"00328DA9", x"002F7896", x"FF2414CD", x"00502C13", x"FF1322C1", x"FFE8137B", x"FF32D64E", x"FF068968", x"FED786C0", x"FEC38C6C", x"FE856C80", x"FE81C28A", x"FEAE8310", x"FE12B1B8", x"001D7ACE", x"FFACDEB2", x"FE4618A0", x"FE69CD04", x"FF1F1F23", x"003FA8DC", x"00EE6DF9", x"FFC3C9C5", x"00A652F5", x"FF5FB213", x"FFC33900", x"FFD29B78", x"FEE327DA", x"000186C0", x"004D6F0E", x"00B25345", x"FF1D8EF0", x"FFA71085", x"0009471D", x"0019403F", x"00256FEE", x"FF118093", x"00C5BC7A", x"FECCA736", x"FF651D3C", x"005778E1", x"FF79B0E3", x"FF38FB1A", x"FEAC160A", x"00981435", x"FFCBC3C2", x"006AE687", x"00160792", x"FF1540A6", x"FF8F959E", x"00CDF76E", x"FF703BF9", x"FF791AA9", x"00A06C75", x"FF81331E", x"002FC2B4", x"FF71C47B", x"005A0EF0", x"001DC302", x"FF17C4E6", x"FF22170B", x"006B69D9", x"FF9FB7FB", x"009F8F4B", x"000E17E7", x"FF9A71C7", x"FFCAD755", x"FF781671", x"008BA808", x"00E1C62B", x"FFEEF5A2", x"FF3D1120", x"00CBC8A7", x"00E752B8", x"00C2B54A", x"FFF7D56B", x"004652D6", x"000DE6C5", x"FF8FE4C0", x"FEDE3BF0", x"FFDC3D49", x"007E89C9", x"00AAA91C", x"004595C2"
--  0.032396, 0.005525, 0.004403, 0.002548, -0.012557, -0.009343, 0.002370, 0.026884, -0.010066, -0.009346, 0.006799, -0.013072, 0.031310, 0.027157, 0.001439, -0.023098, 0.009995, 0.030288, 0.011766, 0.014970, -0.018904, -0.035182, -0.013430, 0.001141, 0.031731, 0.007457, -0.006547, -0.008974, -0.006829, -0.019205, -0.014952, 0.006635, 0.024196, 0.030369, 0.014445, -0.022864, 0.035638, 0.037981, -0.005563, 0.008101, 0.040560, -0.006379, 0.020886, 0.009619, 0.023353, 0.016277, 0.038563, 0.032549, -0.022550, 0.022550, -0.006524, -0.018508, 0.005990, -0.004861, -0.023274, -0.031524, -0.019904, 0.003677, 0.021767, 0.021043, 0.009952, 0.034031, -0.029008, -0.016925, 0.025471, -0.015147, 0.064072, 0.044797, 0.037369, 0.089441, 0.078678, 0.089426, 0.085432, 0.051243, 0.085411, 0.049129, 0.033695, 0.032690, -0.015735, -0.016623, 0.034951, -0.023349, 0.019298, 0.021585, -0.028995, -0.004093, -0.000386, 0.026581, -0.009398, 0.032707, -0.026686, 0.022939, 0.034680, 0.012900, 0.029851, 0.030520, 0.072763, 0.092710, 0.091155, 0.151581, 0.134952, 0.150992, 0.181172, 0.147133, 0.124705, 0.092744, 0.017053, 0.019797, 0.040669, -0.020990, 0.004980, 0.026530, 0.003943, -0.008008, 0.012893, -0.029589, 0.029396, 0.027126, -0.010615, -0.011932, 0.001255, 0.050431, 0.008447, 0.024389, -0.019341, 0.036252, 0.061336, 0.074869, 0.102267, 0.146304, 0.189151, 0.164929, 0.108433, 0.052990, 0.073896, 0.010261, 0.030773, -0.005520, 0.000487, -0.027986, -0.013606, 0.002947, -0.034494, -0.007988, 0.019635, 0.019215, 0.016344, -0.022943, -0.001358, -0.032693, 0.009702, -0.025197, -0.003515, -0.046858, 0.000163, 0.003154, 0.049265, 0.050378, 0.042627, 0.038946, 0.010147, 0.030421, -0.017656, -0.008119, 0.018854, 0.031937, -0.009061, 0.024979, -0.002706, -0.007147, -0.004302, -0.018033, 0.005329, -0.011064, -0.036440, 0.003834, -0.035036, -0.046102, -0.026379, -0.053796, -0.077252, -0.106945, -0.092841, -0.091989, -0.035209, -0.060259, -0.042870, -0.044595, -0.058688, -0.059493, -0.059637, -0.022204, -0.048788, -0.024750, 0.026650, -0.006824, 0.028812, 0.021139, -0.007718, -0.031775, 0.021239, -0.013898, 0.006243, -0.056939, -0.020405, -0.062462, -0.056286, -0.094023, -0.111614, -0.097554, -0.057555, -0.081507, -0.120250, -0.118451, -0.172840, -0.190008, -0.122775, -0.090081, -0.054756, -0.030410, 0.002509, -0.027682, 0.001981, -0.013047, -0.004757, 0.028209, -0.028831, 0.015537, -0.031035, -0.023212, -0.037522, -0.044241, -0.024104, -0.050731, -0.024056, -0.074293, -0.056499, -0.087305, -0.096567, -0.074485, -0.175658, -0.238432, -0.248652, -0.229080, -0.175752, -0.154382, -0.117465, -0.051179, -0.024883, 0.012763, -0.000420, -0.009583, -0.007644, -0.007365, -0.012232, -0.017520, -0.022943, -0.015033, -0.015544, 0.007317, -0.046947, -0.002994, -0.046006, -0.081259, -0.018193, -0.045777, -0.051882, -0.106978, -0.198794, -0.235590, -0.287273, -0.210273, -0.163173, -0.114504, -0.110087, -0.053980, -0.025798, 0.015236, -0.026280, -0.033160, -0.032352, 0.004581, -0.028335, -0.011976, -0.030335, -0.016279, -0.044635, 0.018961, -0.031429, -0.032280, -0.007870, -0.049753, 0.015269, 0.012114, -0.061564, -0.125598, -0.228144, -0.220672, -0.224792, -0.165259, -0.102422, -0.051713, -0.071218, -0.061103, -0.043678, -0.003041, 0.010492, 0.018285, 0.015490, 0.034521, -0.027878, -0.033017, -0.023685, 0.012960, -0.032718, 0.040195, 0.023083, 0.036129, 0.042083, 0.055360, 0.091629, 0.025951, -0.094581, -0.155765, -0.137664, -0.148806, -0.135908, -0.104630, -0.067548, 0.014486, -0.010555, 0.058674, 0.004691, -0.026710, -0.015717, -0.022107, -0.031037, 0.003459, -0.008668, -0.020270, -0.019192, -0.016304, 0.023208, -0.002732, 0.030924, 0.028715, 0.002224, 0.100582, 0.063131, 0.029619, -0.080669, -0.122975, -0.054604, -0.091045, -0.058839, -0.061809, -0.007083, 0.072895, 0.107448, 0.052351, 0.020531, -0.019265, -0.005755, -0.029845, -0.028269, -0.007895, 0.034025, 0.002734, -0.028132, 0.016048, 0.041645, 0.056271, 0.045029, 0.045922, 0.095747, 0.116869, 0.088558, -0.009624, -0.083637, 0.001317, 0.012563, 0.032163, 0.019118, 0.036547, 0.070636, 0.122451, 0.096961, 0.089529, 0.046947, -0.014567, 0.023073, 0.002786, -0.009053, -0.016032, -0.031921, -0.000211, 0.015267, 0.012621, 0.043878, 0.065576, 0.071440, 0.078941, 0.081830, 0.140047, 0.014283, -0.058289, 0.004634, 0.070282, 0.048794, 0.039489, -0.044224, 0.021804, 0.077992, 0.114436, 0.104772, 0.079841, 0.082958, 0.013606, -0.019797, 0.034314, -0.007458, -0.006609, 0.009049, 0.025399, -0.036346, -0.018494, -0.003381, 0.029129, 0.064467, 0.110009, 0.163125, 0.097525, 0.056385, 0.029925, 0.048092, 0.069325, 0.051241, -0.033377, 0.012762, 0.010677, 0.071069, 0.130239, 0.127819, 0.067387, 0.014873, -0.030793, -0.035985, -0.007967, -0.027728, -0.003614, -0.019281, 0.014256, -0.000360, 0.001177, -0.024838, 0.021747, 0.099543, 0.134905, 0.206654, 0.117568, 0.084773, 0.008041, 0.018384, 0.014698, -0.044791, -0.062701, 0.021726, 0.071221, 0.099121, 0.098210, 0.083595, 0.034673, 0.054171, -0.024207, -0.037528, 0.029577, -0.002880, 0.023983, -0.012494, 0.019823, -0.056523, -0.022963, 0.001722, 0.037571, 0.125998, 0.168678, 0.189375, 0.205090, 0.068327, 0.047218, -0.017084, -0.052724, -0.064517, -0.023371, 0.022193, 0.076439, 0.064360, 0.058109, 0.026645, 0.004013, -0.012536, 0.021195, -0.030167, -0.027634, -0.029077, 0.033400, -0.005240, -0.019683, -0.015656, -0.080460, -0.060229, 0.043782, 0.111933, 0.150350, 0.238674, 0.235592, 0.166950, 0.049359, 0.034524, -0.004025, -0.004034, 0.091965, 0.090778, 0.118356, 0.058748, 0.058934, 0.019304, -0.035409, -0.029631, -0.009918, -0.023149, 0.004407, 0.018859, 0.004151, -0.036020, -0.010859, -0.051985, -0.054908, -0.095856, -0.052847, 0.041273, 0.157245, 0.227734, 0.263464, 0.208512, 0.094968, 0.076053, 0.092179, 0.134295, 0.163561, 0.146090, 0.120279, 0.059710, 0.010855, 0.021044, 0.003238, -0.002716, 0.014538, 0.014302, 0.031166, 0.031068, -0.029135, -0.034617, -0.027832, -0.004898, -0.030841, -0.080685, -0.093992, -0.043031, 0.071375, 0.196141, 0.242013, 0.225516, 0.251485, 0.230242, 0.175110, 0.156454, 0.158066, 0.072009, 0.075458, -0.000328, -0.025957, -0.055131, -0.063628, -0.009346, -0.018965, -0.022015, 0.028468, 0.006622, -0.009584, -0.033598, -0.025854, -0.033978, -0.035834, -0.113617, -0.071570, -0.048524, -0.032247, -0.002684, 0.121963, 0.168035, 0.214698, 0.185337, 0.161237, 0.088294, 0.052652, 0.019893, -0.054672, -0.038364, -0.012896, -0.006943, -0.016887, -0.015920, 0.011555, -0.031774, -0.010757, 0.030977, 0.004596, -0.000773, -0.030837, -0.034222, -0.024399, -0.084734, -0.097026, -0.128389, -0.113866, -0.107880, -0.126710, -0.047233, -0.045896, -0.065796, -0.031848, -0.095078, -0.111063, -0.074006, -0.085105, -0.064117, -0.065280, -0.031546, 0.015807, -0.037440, -0.025563, -0.007931, -0.028265, 0.006685, -0.007097, 0.026937, -0.036446, -0.002739, 0.004340, -0.021030, -0.059359, -0.047367, -0.141429, -0.116242, -0.165657, -0.169305, -0.156584, -0.167848, -0.147320, -0.133699, -0.132967, -0.055000, -0.020537, -0.017365, -0.026048, -0.043294, -0.006643, 0.006737, -0.028558, 0.030307, -0.000940, 0.009754, 0.031507, 0.015498, -0.019469, 0.012213, 0.017559, 0.009186, -0.034638, -0.028352, -0.074345, -0.070868, -0.108209, -0.071516, -0.059743, -0.123889, -0.093805, -0.077655, -0.073960, -0.003590, -0.052952, -0.035195, -0.039581, -0.005491, -0.028998, -0.024836, 0.035413, 0.015951, 0.015152, 0.025328, 0.006171, 0.005795, -0.026846, 0.009787, -0.028914, -0.002920, -0.025044, -0.030452, -0.036191, -0.038629, -0.046213, -0.046660, -0.041197, -0.060218, 0.003599, -0.010148, -0.053943, -0.049585, -0.027451, 0.007771, 0.029105, -0.007350, 0.020303, -0.019568, -0.007419, -0.005541, -0.034771, 0.000186, 0.009452, 0.021768, -0.027642, -0.010856, 0.001133, 0.003082, 0.004570, -0.029113, 0.024138, -0.037518, -0.018907, 0.010678, -0.016395, -0.024294, -0.041493, 0.018564, -0.006376, 0.013049, 0.002689, -0.028656, -0.013723, 0.025142, -0.017550, -0.016467, 0.019583, -0.015479, 0.005830, -0.017362, 0.010993, 0.003633, -0.028348, -0.027089, 0.013112, -0.011753, 0.019478, 0.001720, -0.012397, -0.006489, -0.016591, 0.017048, 0.027560, -0.002080, -0.023796, 0.024876, 0.028238, 0.023768, -0.000997, 0.008584, 0.001697, -0.013685, -0.035372, -0.004365, 0.015447, 0.020833, 0.008494
--  Sum of weights (converted): FFFFFFFFF72FCACE
    );

    constant weights_n7 : weight_array := (
     x"00856A17", x"00B72313", x"FFC77057", x"00BF0C6E", x"FFF9DAD0", x"FF986287", x"FF8E6324", x"FF557D0B", x"FF1EA976", x"004305C9", x"010E59DE", x"00299759", x"00278391", x"FF91CE87", x"FF8C4081", x"FFA448A7", x"00654515", x"003270F2", x"FF948117", x"003953F4", x"FFCCE20C", x"FFEC123A", x"00CF73C7", x"FF861607", x"0110FC70", x"FF5FF919", x"010F0EAA", x"006DE977", x"007579D7", x"FFBD1319", x"FFB044B9", x"FF29FE94", x"FEE76D9C", x"00CCD619", x"011B5506", x"0052720F", x"FF8BE4F4", x"003DD88B", x"FFF29BA1", x"FEFF3FEA", x"FF10AA9E", x"0062051D", x"FFA78C72", x"FFB76048", x"FF4C4B80", x"007E9722", x"FF6B3B1E", x"FFA20355", x"009C223C", x"01192260", x"0104BF3C", x"007322A6", x"000A6496", x"00DBE41E", x"0102ACE8", x"00835903", x"00560112", x"00468C92", x"001DC578", x"00C10AEE", x"00527B35", x"FF093EF7", x"FF5228DC", x"FEF2E2C8", x"FFA203AB", x"0004623E", x"FF72C665", x"FEDC7300", x"FF258930", x"005CF6BB", x"FFC941D7", x"FFADF6BC", x"00105DCE", x"FFA6D12E", x"FF4B55B0", x"FF6B3966", x"FF80F4B7", x"FEEA219C", x"FEEFD21E", x"FF906E2C", x"006D8FB5", x"011E197E", x"FFF814CE", x"00C7CBEC", x"0060BD82", x"FF16FB9F", x"FF6DA147", x"FFAF8521", x"FF0E6C98", x"0027A783", x"004130F9", x"FF0E4598", x"FFA68930", x"FED35570", x"00E2A123", x"00571390", x"FF2F8EDA", x"0085EB74", x"FEC88CA6", x"006E1F65", x"FF0EDAA0", x"FFE843C1", x"0079539D", x"004CF628", x"001F790A", x"FFC5C6C4", x"FFF66662", x"00F3EECC", x"FF9E5675", x"FFA0F5D5", x"00255836", x"FF720B09", x"FF9162D2", x"0016DC89", x"00DC08CB", x"005F932A", x"FF49A0F4", x"00A5B7E1", x"FF7EE5A0", x"00192453", x"FFB4E401", x"00393361", x"FEE0A680", x"FE5F7F22", x"FE37738C", x"FE195F3A", x"FD56224C", x"FE9ABA34", x"FD5E72B0", x"FE7CB1A4", x"FDC9D0EC", x"FEDE6746", x"FF0B4953", x"FF121155", x"00505FF6", x"FED8C27C", x"0011465C", x"FFE0F2A2", x"FF666CB5", x"00E37B46", x"00B7AA91", x"0058698B", x"0005A04D", x"00A19973", x"FF79BB33", x"FF04B949", x"00E73F82", x"FF2DD9CD", x"FF988A96", x"FEF81DCA", x"FF4C19AC", x"FEAAA394", x"FBD9FB00", x"FBB30C10", x"FA45F038", x"FBC44F78", x"FC4C92B0", x"FB3C5B38", x"FC981840", x"FCE3D254", x"FD98290C", x"FF763363", x"FE028C8C", x"FF47A9F3", x"FFBEBAF8", x"FEEA7D42", x"0072E00D", x"00C2ED26", x"FF1797EF", x"007131CC", x"FFF30D4F", x"0120FFD8", x"FEFA04A0", x"011FA6F4", x"FFCFA4C0", x"01322DB6", x"FFC7AB59", x"004C2552", x"0005178E", x"FF9CFD41", x"FE08513A", x"FCA1AA94", x"FAD00208", x"F9BE52C8", x"FAE18878", x"FC491A70", x"FCA7D7BC", x"FBEA8E70", x"FE2F957C", x"FEC50DC4", x"FE7564F0", x"FF986E9F", x"FF5C360B", x"FFE0F2E4", x"FF2CE1D6", x"FFDA3EE4", x"011E6C30", x"00B68270", x"FF286B15", x"0039DF7D", x"0148217A", x"0098C1AB", x"01AD0B4A", x"02F8C674", x"03C5AB68", x"04234CC0", x"02498580", x"01477074", x"01E894F6", x"FFA60BFE", x"FFCF2603", x"FFAC0D61", x"FF39287D", x"008EBE0C", x"0089B49B", x"FF7C48D1", x"009D43B8", x"FF481A7D", x"FEC14500", x"FE0114DE", x"00102CC8", x"FE6A62AE", x"00C0F91D", x"FF9801F1", x"FFC9E4DF", x"003506EA", x"017866C6", x"001B696C", x"0083BCA9", x"02D7ECAC", x"029D88D8", x"03CB9038", x"05561870", x"04702B98", x"05A4EC30", x"042E5F20", x"04DFB5E0", x"048E2C10", x"0410CD78", x"047E48F0", x"065E1758", x"05FC8508", x"045F3ED8", x"03F94C34", x"01742EA2", x"00CC65EE", x"FF75BE95", x"FF224195", x"FF0CB8B2", x"FF884360", x"005BB071", x"00D9CF4D", x"00B6EBE1", x"FF9E585E", x"01889DF4", x"0208B300", x"0260DCB0", x"02CFE898", x"02BD5468", x"035109EC", x"0435BA00", x"036156FC", x"04AA1760", x"03296964", x"0344A0C8", x"04434D10", x"06B40430", x"08589180", x"07B61D50", x"078918B0", x"06AF6660", x"047FC6D8", x"01C70B74", x"01B59014", x"FF72404D", x"FF8D8956", x"FFB7EBBC", x"00A2426E", x"FEF07AEA", x"00DCFD00", x"002E344A", x"011F508A", x"01B0C788", x"0108CAC2", x"01F3C41C", x"026B3ED4", x"03C968F8", x"0265FDFC", x"03298CF4", x"02E60DF0", x"03690978", x"02EC6C00", x"03469F3C", x"0296D5D4", x"03CC0440", x"04F665C0", x"085A7650", x"07F1CFB8", x"06A87B80", x"053C3A98", x"03226998", x"02574360", x"0021DBAC", x"005E28CF", x"FE7BE200", x"FEB51C7E", x"0055DF9A", x"0112B2FC", x"FF97B8EC", x"0135ED16", x"002ED31D", x"005ECB04", x"01C27C44", x"02A4CA14", x"0146CD72", x"02B01418", x"009B49A6", x"00490D27", x"FFA41407", x"FEACF9C6", x"00B3C1BF", x"FF761505", x"FFDE97CB", x"01BD1B56", x"05C6C638", x"0638E708", x"05BC1538", x"0395635C", x"03486A6C", x"01C90848", x"016D7186", x"FFE08291", x"00757164", x"00A6A60A", x"00283B6B", x"FEE72354", x"003C91AB", x"FF3BF6DC", x"00A1A07F", x"00E12584", x"0268A15C", x"0093CA51", x"FFD280CC", x"00FC9F30", x"00B70D7A", x"FE59DBC0", x"FD386E08", x"FCA6DE6C", x"FB4891D0", x"FA6CF450", x"FBEB4E28", x"FF765879", x"024A21A4", x"04B86028", x"03E9BEF0", x"029836E4", x"01D5D054", x"FFA3E1A5", x"0091AFA6", x"FEEDCAE0", x"FEB350D0", x"FFD11FC4", x"FF890314", x"FF474CFF", x"FFC2662A", x"FFEC5AF5", x"0098749D", x"00C6C43C", x"00C47968", x"00D9BFAF", x"FF2CCADD", x"003E52A6", x"FED66EF8", x"FD1736FC", x"F9326A90", x"F916E738", x"F7722280", x"F58079F0", x"F93C6AC8", x"FCBC8C58", x"017C376E", x"03A51278", x"037E9294", x"03603D48", x"007D2B56", x"01A2EDE8", x"0020677B", x"FFA057F9", x"FEDD9DC8", x"FF654E53", x"011AE6AC", x"00D8B99D", x"00E40963", x"FFEC11ED", x"FF7BD068", x"009468BC", x"FFE6A93C", x"FF6836B9", x"FFACC3B5", x"FF3F8FFB", x"FC22BED8", x"F9C04990", x"F8B25E38", x"F68C5120", x"F5635C30", x"F57A4BF0", x"F8682E70", x"FD65743C", x"028AD24C", x"03BBA610", x"03DFEDDC", x"02BD5494", x"01AAC25A", x"019CFB0A", x"006C27E5", x"FED534FE", x"FFF2313E", x"009EC8D9", x"FFB30A19", x"FFC95BD1", x"FFD85E70", x"00B3AC13", x"00FA0FFB", x"FF42E2DF", x"00E1EA65", x"0020918E", x"FF6D5ACE", x"FD35C8B0", x"FB9330C8", x"FBB69DE8", x"F9706CB0", x"F800F428", x"F76FEA70", x"F8E5D178", x"FB2C5E90", x"00E49B7B", x"0277BC04", x"04613D40", x"044C9D28", x"0259F0CC", x"01DA699E", x"01570514", x"FF535E74", x"FFADD1FB", x"FFF485B4", x"00E5F738", x"003D8CBC", x"FF06EDCD", x"FFAAA4F4", x"01210A98", x"FFD90805", x"00E8A9F6", x"0027E2A3", x"002E8030", x"FE4C7C84", x"FEEF2CBE", x"FCC807D0", x"FB450440", x"FB7F3DC8", x"FAB75850", x"F9DA0648", x"FBEDC088", x"FFED28AE", x"028DD7C8", x"02F3C1F8", x"02AC6710", x"01B9BDFC", x"021C9CC8", x"0103F2EE", x"FF1FD42C", x"FF6F132F", x"FFD190DB", x"FEB4041A", x"00DE6AF5", x"FFDCC0D3", x"FF88D9D9", x"002093B7", x"0069A649", x"003CC5D8", x"010A8A2A", x"007DE196", x"FF24C901", x"FE8FBD46", x"FDCCDA84", x"FC615780", x"FB384348", x"FB63A870", x"FB614000", x"FBFD1F90", x"FFEDB317", x"0191D478", x"040A7F40", x"02811480", x"01BEF350", x"008A36D3", x"FFA96E6F", x"FF826F90", x"FF95B185", x"FECED20A", x"FED97E50", x"FFEA060E", x"FF631324", x"FFF12E92", x"0054F6FE", x"00833D16", x"FEE4F960", x"006E8E32", x"FF78F8E1", x"FEDA46E0", x"FE63DA92", x"FDD29FC0", x"FDBD82FC", x"FB9CD1D8", x"FC680780", x"FCDDCC8C", x"FC2F9DB0", x"FF233AB1", x"01394AE6", x"03310AA8", x"02835A30", x"FFA22A4C", x"FF699623", x"FF4674F9", x"FDB41CB0", x"FCD2A260", x"FDEEAEC0", x"FEA19896", x"FF431CD2", x"FF694DC3", x"FFA1FB49", x"FF6EF2F5", x"00BCE597", x"FF5AB9D7", x"FF9ECD22", x"00BE1D00", x"FF530D26", x"FF644E40", x"FE3434C8", x"FCAFD50C", x"FD7A8C70", x"FBD68FF8", x"FB7A6D68", x"FC1EB1D8", x"FE1B5B7C", x"01315754", x"030AED90", x"02550394", x"FFA53F34", x"FECCF77C", x"FDABCA00", x"FDC86D84", x"FC7D6D90", x"FBD7EE10", x"FDDA3588", x"FDFA7454", x"FF617D0F", x"FFF7AB91", x"00505A28", x"009F3718", x"FF32D4AE", x"FF11B0E2", x"01122042", x"0101D7FE", x"FF5B3E74", x"0080E5E9", x"FEE7D5D4", x"FD5D3BB4", x"FC30641C", x"FBB063B0", x"FD1C97CC", x"FC5F62AC", x"FE2062EC", x"01C3EC0C", x"00DD3F2A", x"01E4E854", x"FFDA170D", x"FE6DC34E", x"FD517CDC", x"FC1BBAA8", x"FCE5E444", x"FD2FC94C", x"FD10F478", x"FD8CCB1C", x"FE3F4604", x"FF959600", x"00450024", x"FF4463E9", x"0035E5F1", x"00A8887F", x"00ABEE65", x"FF88E8AE", x"0011F343", x"FE7AAC6E", x"FFC16F79", x"FD34C8DC", x"FD687374", x"FCA3ABB4", x"FC3E04A0", x"FCFB915C", x"FE9277A6", x"FF5B8503", x"00DA5DBA", x"FF4256E7", x"FE15FAD4", x"FE0B4F7A", x"FCD3E53C", x"FC8852B4", x"FDB20488", x"FC5DB5E0", x"FD3B1D78", x"FF282BF5", x"0031B08C", x"FEB62842", x"0051C120", x"01206534", x"FFD0FEF0", x"FF535C12", x"008F85E0", x"009D2B52", x"FFBE95EC", x"FEC55550", x"FF8EFEA8", x"FE4FA26C", x"FDC487AC", x"FF46E0CA", x"FF81F203", x"FFA6A6D2", x"FE89470A", x"0079A1D2", x"00092DA5", x"007D1FAF", x"FF5BEAE7", x"FEB607B4", x"FD3EE76C", x"FE65BC96", x"FD800E6C", x"FCECE208", x"FFCD22F5", x"FF16D094", x"00480955", x"FFB1C2E1", x"FFC7A8F0", x"0100FCA6", x"00F2EA66", x"FF777334", x"00092419", x"00C19F56", x"FFFED038", x"FFD470F7", x"01278BC2", x"014525DA", x"0032707F", x"01362606", x"007C1A9B", x"00E1A8FE", x"017E411C", x"001C0892", x"001E4D72", x"00963D15", x"FFC2F99E", x"0134C91A", x"FECA9B28", x"FDEB51B8", x"FE9A6A20", x"FE93D95C", x"FF1EBD78", x"FF8E25D9", x"00D4647E", x"FECB36A4", x"FF45D2AF", x"00359D1E", x"FEFB8AC6", x"FF18DC38", x"00E02E8C", x"0070356E", x"FFAC3ABB", x"008DBB0E", x"00D551E7", x"010725E8", x"02D5B3C8", x"026963CC", x"039269E8", x"023624B4", x"026DBDC4", x"02E70A84", x"039AAF80", x"02A6FD70", x"03B038FC", x"013C2C34", x"00BA5BFB", x"00C3E213", x"FE7F3D04", x"FE3A6E36", x"FF31A6F9", x"FEAE9FAA", x"0014B966", x"FFB6C3DC", x"FFA11B5C", x"00A1C5EA", x"00110599", x"FEF83AC4", x"FEEAC146", x"00B72A7B", x"008827A9", x"00D4BB68", x"FF868AAE", x"00D87B1D", x"02FD1CC0", x"03F01F98", x"0464B3B8", x"050C2D50", x"04136908", x"03A2673C", x"0532C9A0", x"053EC120", x"03CD64A4", x"0311EDE8", x"01F7EC70", x"FFC794E4", x"FF8B02F4", x"FF54200D", x"00383D99", x"FF89AE2F", x"006AB0C2", x"0103BF54", x"FFC14386", x"FFB8AC61", x"FF483C7B", x"FFE9ABEE", x"FEF44258", x"00C5C1D7", x"00FC4A3A", x"0052B3DA", x"012D582C", x"00E5EBEB", x"01818AA8", x"025A85D0", x"00F58646", x"0231F31C", x"031CBE24", x"02773628", x"02314894", x"028BFEDC", x"022EFE98", x"01EC15B4", x"00CDCAF2", x"009F4AE2", x"00F5F85C", x"FF69B266", x"007932D4", x"FF194311", x"FF47A05E", x"001E40E5", x"010F5D2C", x"FEF1CE38", x"007F5970", x"00332B60", x"FF10F02B", x"FF2B92B9", x"009367C3", x"FF6E1934", x"00D1353B", x"FF3F3A8F", x"00EC3C98", x"FF840AB4", x"00997BB2", x"0089DF86", x"FF53E832", x"FFC0679E", x"003DD8E8", x"00A6CB03", x"01250FA8", x"001D897F", x"00B80C24", x"FFBC9156", x"FF993370", x"00C65483", x"FFB55D48", x"FF0B3D91", x"000E7D95", x"FFD64AD9", x"00532CA2", x"FF6AC0D2", x"000C99F9"
--  0.016286, 0.022356, -0.006904, 0.023321, -0.000750, -0.012648, -0.013869, -0.020814, -0.027507, 0.008181, 0.033002, 0.005077, 0.004823, -0.013451, -0.014129, -0.011196, 0.012362, 0.006157, -0.013122, 0.006998, -0.006240, -0.002433, 0.025324, -0.014882, 0.033323, -0.019535, 0.033088, 0.013417, 0.014340, -0.008170, -0.009733, -0.026124, -0.034249, 0.025004, 0.034586, 0.010064, -0.014173, 0.007550, -0.001635, -0.031342, -0.029216, 0.011965, -0.010797, -0.008865, -0.021937, 0.015453, -0.018160, -0.011473, 0.019059, 0.034318, 0.031829, 0.014055, 0.001269, 0.026842, 0.031577, 0.016034, 0.010499, 0.008612, 0.003634, 0.023565, 0.010069, -0.030121, -0.021221, -0.032851, -0.011473, 0.000535, -0.017239, -0.035590, -0.026668, 0.011348, -0.006682, -0.010014, 0.001998, -0.010887, -0.022054, -0.018161, -0.015508, -0.033920, -0.033225, -0.013619, 0.013374, 0.034924, -0.000967, 0.024389, 0.011809, -0.028444, -0.017867, -0.009824, -0.029489, 0.004841, 0.007958, -0.029508, -0.010921, -0.036702, 0.027665, 0.010629, -0.025445, 0.016348, -0.038019, 0.013443, -0.029437, -0.002897, 0.014810, 0.009395, 0.003842, -0.007107, -0.001172, 0.029777, -0.011922, -0.011602, 0.004559, -0.017329, -0.013503, 0.002791, 0.026860, 0.011667, -0.022262, 0.020229, -0.015760, 0.003069, -0.009169, 0.006983, -0.035077, -0.050843, -0.055731, -0.059403, -0.083236, -0.043612, -0.082221, -0.047279, -0.069114, -0.035351, -0.029872, -0.029044, 0.009811, -0.036040, 0.002109, -0.003791, -0.018747, 0.027769, 0.022420, 0.010793, 0.000687, 0.019726, -0.016390, -0.030673, 0.028229, -0.025653, -0.012629, -0.032212, -0.021960, -0.041670, -0.129641, -0.134394, -0.178963, -0.132286, -0.115653, -0.148882, -0.106434, -0.097190, -0.075176, -0.016821, -0.062189, -0.022502, -0.007967, -0.033876, 0.014023, 0.023795, -0.028370, 0.013818, -0.001581, 0.035278, -0.031980, 0.035114, -0.005903, 0.037375, -0.006876, 0.009295, 0.000622, -0.012086, -0.061485, -0.105265, -0.162108, -0.195517, -0.159969, -0.116076, -0.104511, -0.127618, -0.056691, -0.038446, -0.048170, -0.012643, -0.019994, -0.003790, -0.025771, -0.004609, 0.034964, 0.022279, -0.026316, 0.007065, 0.040055, 0.018647, 0.052374, 0.092868, 0.117880, 0.129309, 0.071475, 0.039971, 0.059641, -0.010981, -0.005963, -0.010248, -0.024273, 0.017425, 0.016810, -0.016079, 0.019197, -0.022448, -0.038908, -0.062368, 0.001974, -0.049513, 0.023556, -0.012694, -0.006605, 0.006473, 0.045947, 0.003346, 0.016081, 0.088858, 0.081730, 0.118599, 0.166760, 0.138693, 0.176382, 0.130661, 0.152308, 0.142355, 0.127051, 0.140416, 0.198986, 0.187075, 0.136627, 0.124182, 0.045432, 0.024951, -0.016877, -0.027068, -0.029697, -0.014616, 0.011193, 0.026588, 0.022329, -0.011921, 0.047927, 0.063562, 0.074324, 0.087879, 0.085612, 0.103642, 0.131558, 0.105632, 0.145763, 0.098805, 0.102127, 0.133215, 0.209475, 0.260812, 0.240981, 0.235485, 0.208911, 0.140598, 0.055547, 0.053413, -0.017303, -0.013973, -0.008799, 0.019807, -0.033145, 0.026976, 0.005640, 0.035073, 0.052830, 0.032323, 0.061007, 0.075591, 0.118336, 0.074950, 0.098822, 0.090583, 0.106572, 0.091360, 0.102371, 0.080913, 0.118654, 0.155078, 0.261043, 0.248268, 0.208067, 0.163602, 0.097951, 0.073152, 0.004133, 0.011494, -0.047378, -0.040392, 0.010483, 0.033533, -0.012729, 0.037833, 0.005716, 0.011571, 0.054991, 0.082616, 0.039893, 0.083994, 0.018956, 0.008917, -0.011221, -0.041385, 0.021943, -0.016836, -0.004078, 0.054334, 0.180514, 0.194446, 0.179209, 0.111986, 0.102590, 0.055790, 0.044610, -0.003844, 0.014336, 0.020343, 0.004911, -0.034285, 0.007394, -0.023930, 0.019730, 0.027484, 0.075272, 0.018041, -0.005554, 0.030838, 0.022345, -0.051531, -0.086862, -0.104630, -0.147391, -0.174200, -0.127526, -0.016804, 0.071549, 0.147507, 0.122283, 0.081081, 0.057350, -0.011245, 0.017784, -0.033473, -0.040611, -0.005722, -0.014525, -0.022546, -0.007520, -0.002398, 0.018610, 0.024263, 0.023984, 0.026581, -0.025782, 0.007608, -0.036324, -0.090916, -0.212596, -0.215954, -0.267318, -0.328067, -0.211375, -0.101984, 0.046413, 0.113900, 0.109201, 0.105498, 0.015279, 0.051139, 0.003956, -0.011677, -0.035447, -0.018884, 0.034534, 0.026456, 0.027837, -0.002433, -0.016136, 0.018116, -0.003093, -0.018529, -0.010161, -0.023491, -0.120759, -0.195277, -0.228227, -0.295371, -0.331621, -0.328821, -0.237283, -0.081365, 0.079446, 0.116656, 0.121085, 0.085612, 0.052095, 0.050413, 0.013203, -0.036474, -0.001686, 0.019383, -0.009395, -0.006670, -0.004838, 0.021933, 0.030525, -0.023085, 0.027578, 0.003976, -0.017901, -0.087185, -0.138282, -0.133958, -0.205026, -0.249884, -0.267588, -0.221946, -0.150834, 0.027906, 0.077116, 0.136870, 0.134352, 0.073479, 0.057912, 0.041873, -0.021073, -0.010032, -0.001401, 0.028072, 0.007513, -0.030404, -0.010419, 0.035283, -0.004757, 0.028401, 0.004869, 0.005676, -0.053163, -0.033304, -0.100582, -0.147825, -0.140718, -0.165119, -0.192136, -0.127228, -0.002300, 0.079815, 0.092256, 0.083545, 0.053924, 0.065993, 0.031732, -0.027365, -0.017691, -0.005668, -0.040525, 0.027151, -0.004303, -0.014545, 0.003977, 0.012897, 0.007419, 0.032537, 0.015366, -0.026760, -0.044954, -0.068743, -0.113117, -0.149382, -0.144085, -0.144379, -0.125351, -0.002234, 0.049052, 0.126281, 0.078257, 0.054559, 0.016872, -0.010567, -0.015328, -0.012977, -0.037253, -0.035951, -0.002683, -0.019156, -0.001809, 0.010372, 0.016020, -0.034549, 0.013496, -0.016483, -0.035855, -0.050311, -0.068039, -0.070616, -0.137107, -0.112301, -0.097925, -0.119188, -0.026950, 0.038244, 0.099737, 0.078534, -0.011454, -0.018361, -0.022649, -0.071764, -0.099288, -0.064614, -0.042774, -0.023058, -0.018396, -0.011477, -0.017706, 0.023059, -0.020175, -0.011865, 0.023207, -0.021112, -0.019006, -0.056127, -0.103536, -0.078790, -0.130058, -0.141305, -0.121253, -0.059160, 0.037273, 0.095084, 0.072878, -0.011078, -0.037480, -0.072780, -0.069284, -0.109689, -0.129891, -0.067113, -0.063177, -0.019350, -0.001017, 0.009809, 0.019435, -0.025045, -0.029090, 0.033463, 0.031475, -0.020112, 0.015735, -0.034200, -0.082369, -0.119093, -0.134718, -0.090260, -0.113356, -0.058547, 0.055166, 0.027008, 0.059193, -0.004628, -0.049101, -0.083803, -0.121615, -0.096937, -0.087917, -0.091680, -0.076563, -0.054776, -0.012990, 0.008423, -0.022902, 0.006579, 0.020573, 0.020988, -0.014537, 0.002191, -0.047525, -0.007637, -0.087307, -0.081000, -0.105021, -0.117429, -0.094291, -0.044621, -0.020078, 0.026656, -0.023152, -0.059817, -0.061119, -0.099134, -0.108359, -0.072019, -0.113561, -0.086534, -0.026346, 0.006066, -0.040264, 0.009980, 0.035205, -0.005738, -0.021074, 0.017520, 0.019186, -0.007985, -0.038411, -0.013795, -0.052779, -0.069760, -0.022598, -0.015388, -0.010907, -0.045742, 0.014848, 0.001120, 0.015274, -0.020030, -0.040280, -0.086071, -0.050081, -0.078118, -0.096084, -0.006209, -0.028465, 0.008794, -0.009551, -0.006877, 0.031370, 0.029653, -0.016669, 0.001116, 0.023636, -0.000145, -0.005317, 0.036077, 0.039691, 0.006157, 0.037860, 0.015149, 0.027546, 0.046662, 0.003422, 0.003699, 0.018340, -0.007449, 0.037694, -0.037768, -0.065025, -0.043651, -0.044452, -0.027498, -0.013898, 0.025927, -0.037694, -0.022727, 0.006545, -0.031794, -0.028215, 0.027366, 0.013697, -0.010226, 0.017301, 0.026040, 0.032123, 0.088587, 0.075365, 0.111623, 0.069109, 0.075896, 0.090703, 0.112633, 0.082885, 0.115262, 0.038595, 0.022749, 0.023912, -0.046968, -0.055367, -0.025189, -0.041184, 0.002530, -0.008940, -0.011584, 0.019748, 0.002078, -0.032199, -0.033843, 0.022359, 0.016620, 0.025968, -0.014826, 0.026426, 0.093397, 0.123062, 0.137293, 0.157736, 0.127369, 0.113575, 0.162450, 0.163910, 0.118822, 0.095939, 0.061514, -0.006887, -0.014281, -0.020981, 0.006865, -0.014443, 0.013024, 0.031707, -0.007658, -0.008707, -0.022432, -0.002726, -0.032683, 0.024140, 0.030797, 0.010096, 0.036785, 0.028067, 0.047063, 0.073550, 0.029971, 0.068597, 0.097259, 0.077052, 0.068516, 0.079589, 0.068237, 0.060069, 0.025121, 0.019445, 0.030026, -0.018348, 0.014795, -0.028166, -0.022507, 0.003693, 0.033125, -0.032983, 0.015546, 0.006246, -0.029182, -0.025931, 0.017994, -0.017810, 0.025538, -0.023532, 0.028837, -0.015132, 0.018736, 0.016830, -0.021007, -0.007763, 0.007550, 0.020360, 0.035774, 0.003606, 0.022467, -0.008231, -0.012549, 0.024210, -0.009111, -0.029878, 0.001769, -0.005091, 0.010153, -0.018219, 0.001538
--  Sum of weights (converted): FFFFFFFFDD0CEB1A
    );

    constant weights_n8 : weight_array := (
     x"FF6FA9A2", x"FF4F2E3D", x"0042E139", x"005A6E0E", x"0036203D", x"010E406E", x"001B1F2B", x"0018E11B", x"FFD9C01C", x"FEE52446", x"00726E07", x"00E4132E", x"001CEA07", x"FF1B3DB8", x"01063CA6", x"00418639", x"00D39E71", x"007F11B5", x"002E260B", x"FFA9CC8E", x"003C10C7", x"005E2369", x"FFEE435A", x"FF451F9F", x"FF663DE6", x"FEF3D802", x"FF8D928E", x"FFD0D5A0", x"00EF493C", x"FF637FAB", x"FEE01E1C", x"00A05C47", x"00FC408E", x"FF1BC9D3", x"FFFCED69", x"005C7FA7", x"00BBB46B", x"FFC9E840", x"008348F3", x"00DE3F10", x"00A7CB0A", x"008ABAB4", x"00AD9175", x"FEF5A340", x"003936C7", x"00DDCE1F", x"FF15C28E", x"FEFDE39E", x"FF0D2C82", x"00590AAE", x"010F285E", x"FFE563B5", x"FF8BB214", x"00115080", x"FF0EC3E8", x"0032A582", x"FF3FA62D", x"FF3B13EB", x"FF2A940F", x"FFAD2194", x"00BE5F27", x"003B4F47", x"00CADA91", x"FEE36E56", x"FF0D603E", x"00A928BB", x"00D29A3C", x"00DD2195", x"FEC84014", x"004D3EDC", x"FE9CE030", x"FF63AA9F", x"FFBF5A59", x"0049BABB", x"FF740B56", x"FED88384", x"FECC151E", x"FF7C45FD", x"00D6833D", x"007B79AC", x"008F24F2", x"FF12D5C9", x"FEF91D5C", x"010EB43C", x"00BF1B0A", x"FF81E54B", x"001891D8", x"00D2992C", x"01071280", x"FF129C15", x"FF694942", x"0062B5F7", x"00C36721", x"FFFC2AA7", x"FF92D963", x"FF843AC8", x"0055CA8B", x"FE363F02", x"FF61779C", x"FDEAAEA8", x"FEBC7F74", x"FD91AA10", x"FFA5666C", x"FE7A1E14", x"FF87721C", x"FF010092", x"FFFFD68D", x"FF6CCD02", x"FF666EDA", x"FF800101", x"00B50CFE", x"0028E300", x"FFB4A46E", x"00F92E88", x"00397BF4", x"FFA0E18A", x"FFEF6919", x"FF7C19F8", x"FF61CEC6", x"FF558EAA", x"FFCA7A94", x"FE3E363A", x"FE1E6BBC", x"FF9CF769", x"FE9D949C", x"FF0B4FE0", x"FFE81531", x"FF1E08E4", x"00293E0F", x"FE9F22CC", x"FEA10014", x"FDB098F4", x"FF2AAAA9", x"FE1DB64C", x"FFF03C3B", x"FF6EFB97", x"FF75E9A3", x"FF9E19EA", x"0072D9B6", x"011F147C", x"004F7C97", x"00B35465", x"FF0924FD", x"FFB545DC", x"FF45ACA7", x"FEEEB6F2", x"FFA91867", x"FEC6012E", x"FF188913", x"FE578DB0", x"FDE12DE4", x"FF301534", x"FFBAC881", x"0205AE44", x"0212EFD4", x"04636348", x"041EC370", x"027B1D34", x"01607F66", x"FF8B2BBF", x"008591A7", x"FEE866EA", x"FF09712A", x"FF85A832", x"00450437", x"FFA932F4", x"008D73F2", x"0095E47A", x"FFDBD9C0", x"00C1FA0D", x"FEFE2106", x"FF4EDFDC", x"FFB82C27", x"FF68DB96", x"FF7E4A0A", x"FFAE1EF9", x"FE415520", x"0004CAC5", x"002CFDDD", x"019DBD08", x"01F657E8", x"01A3165E", x"0243829C", x"027AD920", x"034E8AF4", x"0373CF14", x"01C95274", x"01E0D1C2", x"00D3C794", x"00966B18", x"001C43C6", x"FF52AB46", x"FFCFE893", x"00F83E22", x"00F7D60D", x"FF9C0157", x"00F02350", x"00F0441D", x"FF02F924", x"FEC57780", x"FF2D90D7", x"FF54602D", x"FF9F5F94", x"000CFD97", x"00F3FD0A", x"FFFEC144", x"01A97356", x"01017A0C", x"FFAA112A", x"FF44E689", x"FF9F237E", x"009BD916", x"FED05540", x"FF932DC0", x"FF28150E", x"011D6AE6", x"013BFC36", x"0108DF90", x"022B46B4", x"021185FC", x"01863F04", x"001E675B", x"FFFBB641", x"008BE3D8", x"0062A816", x"FF06D64F", x"FF867B3E", x"00983506", x"FF3E2462", x"00ABC0B2", x"FFDF4DD9", x"02012950", x"00D16381", x"030470F0", x"019938B4", x"0203BC08", x"0186E33C", x"00120A2C", x"FDFAA348", x"FDA671C8", x"FCEEEB54", x"FD48DBE0", x"FFB44C4F", x"002B8EFD", x"019508D2", x"02CF8CC0", x"01E720DC", x"024AE7B0", x"01425C78", x"FF37116E", x"00E96D5C", x"001226A9", x"FEEC5CC8", x"FF984BBB", x"00272714", x"00B5CC89", x"FFA33520", x"0148BBAC", x"0082EE13", x"0121370A", x"02DF8658", x"0307C980", x"03B3CC40", x"030DC368", x"0045138C", x"FE81C73A", x"FDA0872C", x"FB3A9BF0", x"FCFC48C4", x"FE313ACA", x"FE5B9026", x"01F25C6A", x"01617BD0", x"03D9B7B0", x"02FD50B8", x"02DDEAE4", x"0254EDCC", x"0055ED7D", x"FF78DFA2", x"00860487", x"FFD07BFE", x"01046A0E", x"FF18E94B", x"FFAC3F3B", x"FF42A2B6", x"FFF9F256", x"0142594C", x"02211C00", x"031945B8", x"0424A298", x"036AD2A4", x"02327448", x"0217D7DC", x"FF3B4DA5", x"FE475AE6", x"FCC70E64", x"FD54F040", x"FE03595C", x"FFE3451C", x"01CD08F2", x"028A6F4C", x"0497DA80", x"045ACFC8", x"038ECCB8", x"01028AE4", x"FF80694F", x"00793BFF", x"0107719E", x"FFD16BB2", x"00EA0B6C", x"00C3A4F1", x"004A5A8F", x"FFD47C71", x"0047CE96", x"01498B64", x"0288682C", x"0351947C", x"02C53AFC", x"0278FB04", x"0287A488", x"0466C050", x"032CC150", x"FF59631B", x"FD6272A8", x"FD51CE54", x"003E9130", x"010EFF4E", x"031C5674", x"02417664", x"04741DB8", x"04004F70", x"0223E6E8", x"00AB5CA3", x"00D35DD9", x"FF86CF0A", x"FF88C08C", x"006DAD56", x"FF1E3E8E", x"00406AD9", x"FFE10701", x"00006AF4", x"0048C29B", x"00C9A134", x"003A848B", x"01A3EA98", x"0052F1B4", x"015475BC", x"0178D410", x"0605F0D8", x"0590B5B8", x"02A62614", x"00A8057C", x"005BE1E1", x"FFB839E8", x"FF839A27", x"0231F36C", x"02D44874", x"020C3538", x"01A1973E", x"00FBACBC", x"00572386", x"00FDB7F6", x"FF63FD09", x"FEEF92E2", x"FFCF9F59", x"FF5506F4", x"FF3B914B", x"FF9ED8BB", x"FFBDA524", x"003A88C7", x"FFC1E0FF", x"FFB22246", x"FF4CF125", x"FE717F5E", x"FE553266", x"01DAB1A4", x"053CAB20", x"064564B8", x"02DA711C", x"01F0632A", x"01E49E9C", x"FFB2FF19", x"FFA454D7", x"FFF25E0C", x"FF5BE535", x"0075F37E", x"FFE96B4E", x"004D60A8", x"0093BCCD", x"FFBD8361", x"00DD33EC", x"000B5017", x"FFC83746", x"00BEF44A", x"00E0D27E", x"FF9D52C5", x"0050B8C2", x"FEBDBCEC", x"FDF43D2C", x"FC409568", x"FBA87F28", x"FBB70E00", x"FCCE68A0", x"018A507E", x"05B82968", x"053654A8", x"04818360", x"033FF450", x"0128AFA2", x"FEFF85D6", x"FC4E77FC", x"FCCE0748", x"FD0F3744", x"FDC03C88", x"FE83EF9A", x"FFD33A0B", x"FE84514C", x"FF54AC36", x"008F62BF", x"00984447", x"FFB523E5", x"FFBC8392", x"FFD4358E", x"00BE6183", x"006DD17D", x"FE29B144", x"FDCFB6EC", x"FBA2F680", x"FB47AD30", x"FC193C4C", x"FDB1BE70", x"0145A944", x"0646DA38", x"0610A170", x"03814C24", x"012F7592", x"FF9A8033", x"FDC033E8", x"FB6CE580", x"FBCFDBD0", x"FCC28448", x"FE05720C", x"FEEF923A", x"FE647596", x"FFEC0B18", x"000ACEA6", x"001BB0CF", x"FF02BBF0", x"010EB6DE", x"0081DCAE", x"001AD7AD", x"00522DCF", x"FF2EF2E2", x"FDBDF2A0", x"FD7B1A40", x"FCA8B4DC", x"FF32D505", x"FFA13F2E", x"015DD294", x"032E7824", x"05781610", x"04E05F98", x"0075CD83", x"0073E25D", x"FFF51373", x"FC2E0010", x"FCB3BA48", x"FB2E86C0", x"FC94A218", x"FE22ACCE", x"FF022811", x"001A6D80", x"006D7944", x"FEA73752", x"001F8BEF", x"FEF95498", x"00A68C63", x"00560AC2", x"00D82E60", x"000F81F7", x"00133D67", x"FE74DC6E", x"FD4D833C", x"FE671F22", x"00F3318C", x"01EACD1C", x"05351AC0", x"0555C818", x"053E25D8", x"03888070", x"FEF8A922", x"FE66AB62", x"FEDC2D74", x"FE12B336", x"FCB46A54", x"FDFF780C", x"FD37A658", x"FE5100F8", x"FD80699C", x"FE3AB6B8", x"FFFF6FDA", x"003DC0BC", x"FF6E590A", x"0065E9D8", x"FFB35801", x"00A331E0", x"00135640", x"FF5FDB29", x"FF38EF10", x"FD8B0808", x"FF766019", x"0171FE50", x"03DA372C", x"042BEB90", x"0529C0F8", x"05062380", x"038D49E4", x"FEF80A06", x"FCFA4D24", x"FDBED694", x"FF195206", x"FE27E9EE", x"FD2EE334", x"FE20591C", x"FE00DD0C", x"FE8ED53E", x"FF3ABF09", x"FEAA58EE", x"FEA90F90", x"FF8194C6", x"00087546", x"00D682E3", x"006A2AC5", x"FF54F51D", x"FEDFA668", x"FFB2972D", x"FEAA1336", x"FF6E3DDB", x"FE6C7A80", x"010BB954", x"024604E0", x"03B772B8", x"0315C224", x"01A0A7AE", x"FFC83439", x"FE3293E2", x"FD73B3E4", x"FE415C5A", x"FE2CDD90", x"FE2CD97C", x"FFFEB7CA", x"FE96A986", x"FE6C7DE0", x"FEB4E64E", x"00878742", x"00CCE07D", x"FF15366E", x"FF066204", x"FEF36454", x"00875B12", x"FF8A2B5B", x"00DA0435", x"FF84E71D", x"006F88E8", x"FF8015FE", x"FF9BD44C", x"00259F78", x"0056542F", x"02077FE4", x"010D8FBE", x"008543DC", x"FFB90466", x"FD808B70", x"FD6DE864", x"FC924384", x"FCCD747C", x"FD14336C", x"FD420CB4", x"FFC2A361", x"FFEDEB78", x"00DA58A0", x"004D343E", x"0052A709", x"FFB2F7ED", x"001DB898", x"FFA91E9F", x"006DF373", x"FF7ADEFE", x"00B8FD87", x"004FFB6A", x"00877A85", x"FF95C25A", x"FF68836F", x"FFFBBBD5", x"FFB6C746", x"015B69BE", x"FFA70D51", x"004FF617", x"FF064902", x"FF9AC666", x"FFBDD7E7", x"FFCEB06F", x"FE97934C", x"FF5653DF", x"FE533DE8", x"FF436948", x"0138B546", x"FF6E809A", x"00A09E6C", x"FF30DFD5", x"0095AE49", x"FEC4921A", x"FE94C802", x"FF91C6B7", x"00E6633D", x"0093D090", x"00BC04FF", x"FFBBD29B", x"00F525A9", x"FF2B6356", x"FF032C8A", x"FDD1A6F0", x"FF3EFD27", x"FFEF72F7", x"FECC98E2", x"00DF5863", x"014CF092", x"03EC4A88", x"03E045A4", x"04B253D0", x"0363575C", x"03483404", x"00EE505B", x"0246F058", x"00E9FBE0", x"01F80BDC", x"FFA722D5", x"FFE14B1C", x"FF8F06EE", x"FF9BF1B5", x"FFCDBA33", x"00535365", x"01059418", x"00AC5732", x"FF72ECBD", x"0112EA08", x"FFD049B5", x"FF35CC74", x"FFC065EB", x"FE87352A", x"FF85F1AA", x"FEC20A5C", x"0046476B", x"007AABF6", x"00F2A694", x"044D5578", x"05D33838", x"07291DE8", x"05F346E0", x"0410C518", x"044C2E20", x"03B3045C", x"00FEF647", x"02096CA8", x"FFFAC552", x"FF4B900C", x"0072510A", x"FFF184C4", x"FF3D5307", x"01018930", x"0016EA0E", x"FF487D8D", x"008636D5", x"0014B52B", x"FFD0A2EE", x"FF1CCF81", x"FF8AF5D5", x"FFCCC019", x"FE360216", x"FF2D3F84", x"FE1430C0", x"FF4D71AE", x"0016676A", x"00824B5A", x"02DB343C", x"0229A700", x"03C9ACE8", x"03256890", x"026AD09C", x"00C385DC", x"00BA2E64", x"011CE8A2", x"01794E1E", x"FF81E5EE", x"FF2F14DE", x"FF75D3EA", x"FF2686F8", x"FFD7A18C", x"FF2F21D1", x"00D4225A", x"00CFA9C5", x"FF45D6C6", x"0101F936", x"00390C94", x"FF2395BC", x"000DE1BF", x"FE6A74EE", x"FE7EAF9C", x"FDDAB2E4", x"FDB7F1D0", x"FDFFC260", x"FE813568", x"FE8BC1D6", x"FD99B970", x"FE1FF32A", x"FF5ACEEC", x"007F24E1", x"0001FE18", x"00BA5AC9", x"FF4F5017", x"0036D832", x"FEE52F0C", x"0087D981", x"FFF1D44D", x"FFE6F305", x"FF61A37A", x"FF001723", x"FF94480B", x"FFE45AC7", x"FF64A114", x"007A491C", x"FFCCFC32", x"00142F1F", x"FEDDF504", x"0033B4B1", x"FF454A1B", x"FEE1C64C", x"FF304DEA", x"FE7E7566", x"FE9BCC94", x"004B15F6", x"006227CE", x"FEB8AE30", x"FFCEAF4E", x"FF04F762", x"00C332BE", x"007FE0F1", x"00539983", x"FEFE48EA", x"FF66B30F", x"FFBFE4B6", x"FEFA37DC", x"FF54F8E8", x"004CF7D0", x"FF11D338", x"004DD817", x"FFF95060", x"FFE7E825", x"FFAA89FE", x"FF62C374", x"FEEE6004", x"FF3873BE", x"00DBFF5B", x"FFE8EDDE", x"011AD1D4", x"000C3CCE", x"FFD74BF4", x"00A986B0", x"FEE43664", x"FF408883", x"009B081C", x"FFA8C3B1", x"00DCC914", x"FFDB01C7", x"00C9DF24", x"000B4E8E", x"001CD5C1", x"FF083713", x"FF9A37AD", x"000E96A8", x"0085AD83", x"0038C497", x"FFC07A5C", x"0001F9AB"
--  -0.017619, -0.021584, 0.008164, 0.011039, 0.006607, 0.032990, 0.003311, 0.003037, -0.004669, -0.034529, 0.013968, 0.027841, 0.003530, -0.027925, 0.032011, 0.007999, 0.025832, 0.015511, 0.005633, -0.010523, 0.007332, 0.011491, -0.002165, -0.022812, -0.018769, -0.032734, -0.013968, -0.005758, 0.029210, -0.019104, -0.035142, 0.019575, 0.030793, -0.027858, -0.000375, 0.011291, 0.022913, -0.006603, 0.016026, 0.027130, 0.020483, 0.016935, 0.021188, -0.032515, 0.006984, 0.027076, -0.028594, -0.031508, -0.029642, 0.010869, 0.033100, -0.003248, -0.014197, 0.002114, -0.029448, 0.006182, -0.023480, -0.024038, -0.026052, -0.010116, 0.023239, 0.007240, 0.024762, -0.034737, -0.029617, 0.020649, 0.025708, 0.026994, -0.038055, 0.009429, -0.043350, -0.019084, -0.007891, 0.009000, -0.017084, -0.036070, -0.037588, -0.016080, 0.026186, 0.015073, 0.017474, -0.028951, -0.032090, 0.033045, 0.023328, -0.015394, 0.002999, 0.025708, 0.032113, -0.028978, -0.018398, 0.012050, 0.023853, -0.000468, -0.013324, -0.015109, 0.010473, -0.055878, -0.019352, -0.065102, -0.039490, -0.075969, -0.011060, -0.047593, -0.014716, -0.031128, -0.000020, -0.017969, -0.018746, -0.015625, 0.022101, 0.004991, -0.009199, 0.030418, 0.007017, -0.011611, -0.002025, -0.016101, -0.019311, -0.020806, -0.006533, -0.054906, -0.058787, -0.012089, -0.043264, -0.029869, -0.002920, -0.027584, 0.005034, -0.043074, -0.042847, -0.072193, -0.026042, -0.058873, -0.001924, -0.017702, -0.016856, -0.011951, 0.014020, 0.035044, 0.009703, 0.021891, -0.030134, -0.009122, -0.022745, -0.033360, -0.010608, -0.038330, -0.028255, -0.051812, -0.066262, -0.025381, -0.008449, 0.063193, 0.064812, 0.137132, 0.128755, 0.077529, 0.043029, -0.014261, 0.016305, -0.034131, -0.030097, -0.014934, 0.008425, -0.010596, 0.017267, 0.018297, -0.004413, 0.023679, -0.031478, -0.021622, -0.008768, -0.018450, -0.015834, -0.009995, -0.054525, 0.000585, 0.005492, 0.050505, 0.061321, 0.051158, 0.070741, 0.077496, 0.103338, 0.107887, 0.055825, 0.058694, 0.025852, 0.018362, 0.003450, -0.021159, -0.005871, 0.030303, 0.030253, -0.012206, 0.029314, 0.029329, -0.030887, -0.038395, -0.025688, -0.020950, -0.011795, 0.001586, 0.029784, -0.000152, 0.051935, 0.031430, -0.010490, -0.022839, -0.011824, 0.019024, -0.037069, -0.013284, -0.026357, 0.034841, 0.038572, 0.032333, 0.067783, 0.064639, 0.047637, 0.003711, -0.000523, 0.017076, 0.012043, -0.030415, -0.014834, 0.018580, -0.023664, 0.020966, -0.003991, 0.062642, 0.025560, 0.094292, 0.049954, 0.062956, 0.047716, 0.002202, -0.063155, -0.073432, -0.095835, -0.084856, -0.009241, 0.005317, 0.049443, 0.087836, 0.059464, 0.071644, 0.039351, -0.024528, 0.028495, 0.002216, -0.033647, -0.012659, 0.004779, 0.022192, -0.011327, 0.040129, 0.015983, 0.035305, 0.089786, 0.094701, 0.115698, 0.095430, 0.008432, -0.046658, -0.074154, -0.149096, -0.094204, -0.056491, -0.051323, 0.060835, 0.043150, 0.120327, 0.093422, 0.089590, 0.072867, 0.010489, -0.016495, 0.016360, -0.005800, 0.031789, -0.028209, -0.010224, -0.023116, -0.000739, 0.039349, 0.066542, 0.096835, 0.129472, 0.106790, 0.068659, 0.065411, -0.024011, -0.053790, -0.100701, -0.083382, -0.062091, -0.003507, 0.056279, 0.079399, 0.143537, 0.136085, 0.111182, 0.031560, -0.015575, 0.014799, 0.032159, -0.005686, 0.028570, 0.023882, 0.009076, -0.005312, 0.008766, 0.040228, 0.079151, 0.103708, 0.086576, 0.077268, 0.079058, 0.137543, 0.099213, -0.020338, -0.081732, -0.083764, 0.007638, 0.033081, 0.097209, 0.070491, 0.139174, 0.125038, 0.066883, 0.020918, 0.025802, -0.014794, -0.014557, 0.013388, -0.027558, 0.007863, -0.003781, 0.000051, 0.008882, 0.024613, 0.007143, 0.051259, 0.010125, 0.041560, 0.046000, 0.188225, 0.173915, 0.082782, 0.020510, 0.011216, -0.008761, -0.015185, 0.068598, 0.088413, 0.063990, 0.050975, 0.030722, 0.010637, 0.030972, -0.019044, -0.033255, -0.005905, -0.020871, -0.023979, -0.011860, -0.008100, 0.007145, -0.007583, -0.009505, -0.021858, -0.048645, -0.052100, 0.057946, 0.163656, 0.195971, 0.089165, 0.060594, 0.059158, -0.009400, -0.011190, -0.001664, -0.020032, 0.014398, -0.002756, 0.009446, 0.018034, -0.008116, 0.027002, 0.001381, -0.006810, 0.023310, 0.027444, -0.012045, 0.009854, -0.039339, -0.063936, -0.117116, -0.135682, -0.133904, -0.099804, 0.048134, 0.178731, 0.162882, 0.140810, 0.101557, 0.036217, -0.031308, -0.115421, -0.099850, -0.091893, -0.070284, -0.046395, -0.005465, -0.046348, -0.020914, 0.017503, 0.018587, -0.009138, -0.008238, -0.005346, 0.023240, 0.013406, -0.057411, -0.068394, -0.136357, -0.147500, -0.121919, -0.072053, 0.039754, 0.196149, 0.189530, 0.109533, 0.037043, -0.012390, -0.070288, -0.142957, -0.130877, -0.101255, -0.061835, -0.033255, -0.050237, -0.002436, 0.001319, 0.003380, -0.030916, 0.033046, 0.015852, 0.003277, 0.010032, -0.025519, -0.070563, -0.078723, -0.104406, -0.025045, -0.011567, 0.042703, 0.099423, 0.170909, 0.152389, 0.014380, 0.014146, -0.001334, -0.119385, -0.103061, -0.150571, -0.106856, -0.058267, -0.030987, 0.003226, 0.013363, -0.042088, 0.003851, -0.032064, 0.020331, 0.010503, 0.026389, 0.001893, 0.002349, -0.048235, -0.084288, -0.049912, 0.029687, 0.059912, 0.162732, 0.166721, 0.163836, 0.110413, -0.032146, -0.049967, -0.035623, -0.060217, -0.102977, -0.062565, -0.086957, -0.052612, -0.078075, -0.055333, -0.000069, 0.007538, -0.017780, 0.012441, -0.009357, 0.019921, 0.002360, -0.019549, -0.024300, -0.076778, -0.016800, 0.045165, 0.120388, 0.130361, 0.161347, 0.156999, 0.110997, -0.032222, -0.094446, -0.070454, -0.028159, -0.057628, -0.088026, -0.058551, -0.062395, -0.045064, -0.024079, -0.041706, -0.041863, -0.015432, 0.001032, 0.026185, 0.012960, -0.020879, -0.035199, -0.009449, -0.041739, -0.017793, -0.049258, 0.032681, 0.071047, 0.116144, 0.096406, 0.050861, -0.006811, -0.056326, -0.079626, -0.054521, -0.057023, -0.057025, -0.000157, -0.044109, -0.049256, -0.040418, 0.016544, 0.025009, -0.028661, -0.030471, -0.032789, 0.016523, -0.014384, 0.026613, -0.015027, 0.013615, -0.015615, -0.012228, 0.004593, 0.010538, 0.063415, 0.032905, 0.016268, -0.008665, -0.078059, -0.080334, -0.107146, -0.099920, -0.091284, -0.085687, -0.007490, -0.002207, 0.026654, 0.009424, 0.010089, -0.009403, 0.003628, -0.010606, 0.013422, -0.016251, 0.022582, 0.009763, 0.016538, -0.012969, -0.018492, -0.000521, -0.008938, 0.042409, -0.010858, 0.009761, -0.030483, -0.012357, -0.008076, -0.006019, -0.043997, -0.020712, -0.052339, -0.023021, 0.038172, -0.017761, 0.019607, -0.025284, 0.018272, -0.038505, -0.044338, -0.013455, 0.028123, 0.018044, 0.022952, -0.008322, 0.029925, -0.025954, -0.030863, -0.068158, -0.023561, -0.002020, -0.037525, 0.027264, 0.040642, 0.122594, 0.121127, 0.146768, 0.105877, 0.102564, 0.029091, 0.071160, 0.028562, 0.061529, -0.010848, -0.003748, -0.013791, -0.012214, -0.006137, 0.010172, 0.031931, 0.021038, -0.017221, 0.033559, -0.005824, -0.024683, -0.007764, -0.045995, -0.014899, -0.038813, 0.008579, 0.014975, 0.029620, 0.134440, 0.182034, 0.223769, 0.185947, 0.127047, 0.134299, 0.115603, 0.031123, 0.063650, -0.000638, -0.022026, 0.013955, -0.001768, -0.023764, 0.031437, 0.002797, -0.022401, 0.016384, 0.002528, -0.005782, -0.027733, -0.014287, -0.006256, -0.055907, -0.025727, -0.060035, -0.021796, 0.002735, 0.015905, 0.089258, 0.067585, 0.118369, 0.098316, 0.075539, 0.023868, 0.022727, 0.034779, 0.046058, -0.015393, -0.025503, -0.016867, -0.026547, -0.004928, -0.025497, 0.025895, 0.025350, -0.022725, 0.031491, 0.006964, -0.026906, 0.001695, -0.049505, -0.047035, -0.067053, -0.071296, -0.062529, -0.046727, -0.045440, -0.074985, -0.058600, -0.020165, 0.015521, 0.000243, 0.022748, -0.021568, 0.006695, -0.034523, 0.016583, -0.001730, -0.003058, -0.019331, -0.031239, -0.013149, -0.003375, -0.018966, 0.014927, -0.006227, 0.002464, -0.035406, 0.006312, -0.022792, -0.034940, -0.025353, -0.047063, -0.043482, 0.009166, 0.011982, -0.039956, -0.006020, -0.030644, 0.023828, 0.015610, 0.010205, -0.031459, -0.018713, -0.007826, -0.031956, -0.020877, 0.009396, -0.029074, 0.009502, -0.000816, -0.002941, -0.010432, -0.019194, -0.033401, -0.024359, 0.026855, -0.002816, 0.034524, 0.001494, -0.004969, 0.020694, -0.034642, -0.023372, 0.018925, -0.010649, 0.026951, -0.004516, 0.024643, 0.001380, 0.003520, -0.030247, -0.012425, 0.001781, 0.016318, 0.006930, -0.007754, 0.000241
--  Sum of weights (converted): 000000005DB9074C
    );

    constant weights_n9 : weight_array := (
     x"00FB80AC", x"00C329EA", x"0063D4B0", x"FF2D2692", x"FF9DA027", x"00BACA25", x"01075DAA", x"FF75AFC9", x"007C50A5", x"FFBB7DE9", x"00B998A7", x"FFD409E0", x"FF17471F", x"FEDD9A9C", x"FFF48803", x"00563B01", x"FF5387E2", x"00E62FFE", x"008AC67C", x"00B06DFA", x"0086CBA5", x"FEE5D162", x"FFCA5B27", x"0097F8F7", x"0090D47E", x"FEF5CC6A", x"FF5A28FB", x"00D54037", x"FF0DC538", x"00DDBD43", x"FFC78D82", x"001576C9", x"008EAEEE", x"004EB930", x"FF43E61F", x"005DCDE0", x"FF02CB44", x"FF698DD9", x"FFC9260E", x"FFBFAEE9", x"00CD02EB", x"FF596D5E", x"00EF2240", x"008149F4", x"0056661A", x"00CA543A", x"FF34C069", x"FF01AE9D", x"00094BC6", x"008F82F5", x"00933C40", x"000C0A59", x"0117D134", x"0067F232", x"007E6B00", x"FF7231B4", x"00593ED5", x"FF927BFE", x"FF13A5F4", x"FF4194EA", x"FF4EFC81", x"FFD3C274", x"FF84803C", x"0108BD4E", x"00729D09", x"FF01A772", x"FFF66435", x"00DC82C7", x"FFC626A3", x"FFF3B646", x"000B5CB2", x"FF5AAA80", x"FEFF9A54", x"FF575AFF", x"FF822651", x"00C02B08", x"FEFD50BA", x"001BB2DF", x"FF89B4B5", x"FFDF00EA", x"FFE57343", x"FF8E48C5", x"004382A7", x"0045253E", x"FF57FD19", x"00B3C2F7", x"0107EA54", x"FF8680C9", x"003B4FB1", x"FF9258F6", x"00C442DB", x"FFDD2650", x"FEE4A0EC", x"001CEE91", x"00AEC439", x"FF9F6D74", x"FF31372F", x"FF49EC73", x"FFD131DE", x"000DC5D7", x"FED0A926", x"FFD218DF", x"0004F0A2", x"008927FD", x"00806862", x"FEDFF1EA", x"FEF97D2E", x"FF043783", x"00B4D15A", x"FF6AF89F", x"00A18085", x"FFD46FF7", x"FF8771DB", x"00DC27D4", x"FFC77BC9", x"FF61CEBA", x"FFD180E4", x"FF3DAD6E", x"FED13B34", x"FFA0740D", x"FF9B5C20", x"FEC5DE54", x"00238F18", x"FE860906", x"FDF88228", x"FEAB93D4", x"FD78C93C", x"FCD24284", x"FD424058", x"FC4B2074", x"FEF3B416", x"FEA3C91A", x"FF347490", x"FE539FBE", x"006407BB", x"FED51F76", x"FF83E7C4", x"FF3E21AB", x"FF6A17ED", x"003E59D4", x"FEDDDA68", x"FEE19450", x"0042CA3A", x"005E8883", x"FFF999AA", x"FF668326", x"FF469F00", x"FF17DC28", x"FE913192", x"FD74ED1C", x"FE8C7CC4", x"FDA69748", x"FBF7D300", x"FBC365C0", x"FA549CA0", x"F9B41878", x"FA4D4CC0", x"F9F16368", x"FAF8AB88", x"FB71DD50", x"FC5A25AC", x"FDA68790", x"FD6B9748", x"FDBE61F8", x"0044F388", x"FFDE09BE", x"00AA90D4", x"00DC0733", x"007FF71E", x"FF9BF83C", x"FFC89973", x"FFE707A5", x"FFE3E30E", x"FF81F5D7", x"FE0986DA", x"FD845D3C", x"FE20A80A", x"FCEA097C", x"FC6A4CE4", x"FE647524", x"FE59EEF0", x"FFFCEEDA", x"030C3B98", x"020A5FA8", x"01984E16", x"016793F0", x"FEF88DEE", x"FD2C9F44", x"FDDECFAC", x"FCE087A4", x"FBFD5918", x"FD066888", x"FE871512", x"FF7F9DEF", x"FF09DEB8", x"FF8F00C7", x"0062E345", x"FEED9412", x"FEE6BB58", x"0026E6AD", x"FFB774DF", x"FDBD0D88", x"FCEE6C2C", x"FDE4A3B8", x"FD997FA0", x"FC276528", x"FEE1020C", x"0093D935", x"03B56970", x"05ACD9A8", x"093101A0", x"0B4E79E0", x"096F1AB0", x"0489A4E0", x"0293A0D0", x"008B81D5", x"FD478524", x"FC0F9B4C", x"FBA53600", x"FC9883A0", x"FDDD5D6C", x"FEA6339A", x"FED3EBB2", x"00B40C61", x"011DA07E", x"00EEDC15", x"009C4FEE", x"0028FAA2", x"FEBCEC08", x"FD8CB6B0", x"FD21A24C", x"FD729924", x"FD802A04", x"FE02F9B2", x"FEFFB634", x"011168D0", x"031DF098", x"0540DE78", x"061531F0", x"06434F98", x"043C96C8", x"0263E208", x"000A585C", x"FFBDE6D6", x"FD8DCEEC", x"FE1EF2DC", x"FC16F3C0", x"FCCCDA34", x"FF7717F9", x"FF0FF12A", x"FFA1CA04", x"0093CA49", x"FF02B69E", x"FFB30572", x"FFCCAACE", x"FFB181D4", x"FEDE3786", x"FDF81FA0", x"FDBD5044", x"FEB12F42", x"003CDC6E", x"00210620", x"02431430", x"03A7F938", x"018204D4", x"02323964", x"0168C46A", x"FF72A210", x"003C58EE", x"006F5DF6", x"00DBF5B1", x"008F6E7F", x"FFB76F19", x"FF47B4F6", x"FD509024", x"FE2F3E7A", x"FFC8412A", x"FF039E20", x"0022FD3C", x"FF66B1B7", x"006AB319", x"0053486F", x"00ABE60C", x"FF94D94D", x"FFE028DB", x"006E6FF5", x"00A6C548", x"00029A3E", x"030391E8", x"023680E0", x"044A9D48", x"024DDD44", x"00D4FBD2", x"FDC5D130", x"FC50AAD4", x"FE29720C", x"FE85661E", x"0002070C", x"015542B0", x"02A63064", x"021F57D8", x"00AA6F5B", x"FFBF6407", x"FF83B1A0", x"FFA0FD34", x"00929CA8", x"0093C33A", x"FF6576FB", x"FFD28E71", x"007CF62E", x"00B83B1B", x"FEBF580C", x"FF5DAFE4", x"00920C6F", x"03477C48", x"0457BA80", x"038155A0", x"03C8923C", x"03CF3498", x"016DCED2", x"FDE3EC18", x"FC4214B8", x"FD57C800", x"FF7BA7DA", x"015DE1EC", x"03AB7B38", x"03D746BC", x"05D78838", x"035B785C", x"01AFFC7C", x"016246B2", x"FF867564", x"FE9C0C9E", x"006E36CF", x"FF7F0916", x"0119F3B8", x"FFAA8A62", x"FF1CFCB1", x"FF063236", x"FFEB81A8", x"0086986D", x"02FC9FB4", x"033ABACC", x"032B9EA4", x"04422038", x"032EA240", x"028EF0A8", x"FFD290DA", x"FCDAEB80", x"FE3692AE", x"00588BC4", x"023188CC", x"03B692CC", x"06657658", x"0609C2B8", x"06C7C638", x"0397A998", x"030AEF20", x"FFCB4729", x"FECFB2E4", x"005F2FCD", x"00C39067", x"FF90B70C", x"00FFEB90", x"0020F07F", x"0066594E", x"FFDB9B5F", x"FFC7A203", x"00BFFB9D", x"0177E578", x"03E45C28", x"0410A6D0", x"04ABE708", x"01EA5F98", x"02183EE0", x"FFD001FD", x"FF891838", x"0059FC50", x"0371AE84", x"04889AF0", x"067889B0", x"0621F5D0", x"07068390", x"05850E68", x"01998AB8", x"01DD9BC4", x"004D1503", x"FE3BE754", x"FE5E0254", x"FFDC1919", x"00E037A9", x"00540F59", x"0028AC20", x"FFEBB169", x"FED4655C", x"00E03E67", x"01D01614", x"00FB8EAA", x"01F7D67E", x"037ECA98", x"023D9498", x"01595F48", x"015770C2", x"0057ACA4", x"0118E2C6", x"0035784A", x"0184C240", x"02C8A120", x"06572A48", x"073AAD60", x"04B4A940", x"019AF1C2", x"FFBA1AE2", x"FE2C0CF0", x"FEE68D92", x"FF88ACE2", x"FE91D4AA", x"FF04F540", x"00D43940", x"002743CE", x"FF75EA1B", x"00BD5D93", x"FF0ABAEB", x"FF9092D1", x"005CE462", x"00DCDB52", x"011AF462", x"01D7C514", x"019B0F14", x"02088958", x"0139B1D2", x"00583957", x"008D6FD2", x"FFA5CD9E", x"FF296381", x"001D7F54", x"05766438", x"04A238B8", x"017F1974", x"FED7D7FA", x"FED21E8E", x"FE4014EA", x"FCAE95C4", x"FE81A190", x"FFB51480", x"0009FC42", x"FFEDD89B", x"FF750E80", x"FF317921", x"FEDF5F54", x"FFF42E6C", x"FF952F1C", x"008C960A", x"FF8DE9BA", x"009862C7", x"FF5FC7FA", x"026732F4", x"018FDACA", x"029CF6FC", x"015946EA", x"00638D32", x"FE6C3B52", x"FE83B536", x"006058A8", x"04AC4458", x"037FD100", x"FEA854E4", x"FDEFDF94", x"FD201EC4", x"FD5B220C", x"FE7BA540", x"FE31C386", x"FE93BE94", x"FF3188BC", x"0017C488", x"FFD43F07", x"FF2E752D", x"0007DD16", x"009EA2B4", x"FFF33B1B", x"00781CE7", x"FEC441F6", x"FFB87E0A", x"FF5FD9D2", x"FF6A7133", x"0103C418", x"016F96B4", x"FFCEBC35", x"FEB27A3C", x"FE29FF1A", x"FDE651B8", x"02687610", x"02839964", x"00190583", x"FE6E3E26", x"FDD70898", x"FDFD89DC", x"FDE2AAA8", x"FCD6E580", x"FD910744", x"FF9AEF4A", x"00DD051F", x"00EF3CDE", x"00726410", x"0115FC28", x"FF798FAF", x"FFED2D58", x"FEDD7896", x"FEBB0910", x"FDE75428", x"FD208174", x"FE208C24", x"FE0F44D8", x"FE547AD4", x"FED0EAF8", x"FCEC8F20", x"FCD2D008", x"FE7F6CB2", x"FF020AFB", x"01CD5212", x"009E503B", x"FE2B5EBC", x"FE400616", x"FE230CE2", x"FE27D1AE", x"FD4CA6F0", x"FE7BD8B4", x"FF6EF187", x"0009F49F", x"FFAF053A", x"FEEED156", x"011E21D6", x"00516B73", x"010216DC", x"0059CEAE", x"FFC26E96", x"FFE6FCBF", x"FF2F0752", x"FD9B3394", x"FD04BC78", x"FBF8B3C0", x"FC0B3F38", x"FB974688", x"FB033D20", x"FCDACA40", x"FE9A9314", x"003562AA", x"FF678B8B", x"FEBD4972", x"FD1F5D88", x"FE9E44E6", x"FDBFCD5C", x"FD926C50", x"FE849856", x"FD75C9E8", x"FF6090AC", x"FF0538EC", x"FFDD7645", x"FF8B7ED2", x"00EC854F", x"FF2689D2", x"00348111", x"FFF78152", x"FEA11E62", x"00319F8D", x"FEE27696", x"FCAEDD1C", x"FB3700D0", x"FBA782A0", x"FB093F90", x"F972C0C0", x"F9D22570", x"FA877160", x"FE564744", x"FDDA9DB0", x"FD536580", x"FDED3020", x"FE34766E", x"FE410C9A", x"FF2D8688", x"FFF0A450", x"FED084C2", x"FF455788", x"FF633005", x"FF247C7E", x"002F7CEB", x"FF64A0EA", x"00A94D8D", x"FF363077", x"FF1079C2", x"FFBD46CC", x"009E1556", x"FE985E9E", x"FE7F69D4", x"FDBE27F8", x"FC0F6578", x"FBF53D58", x"FBAA7840", x"FB0B9A10", x"FA9E44A8", x"FB407A78", x"FC639450", x"FD137050", x"FC5B5C9C", x"FBFCEC28", x"FD659158", x"FD9C188C", x"FF6980B5", x"FEEDC5FA", x"FF775B48", x"FF59A4C2", x"0091948C", x"FEFEC6C6", x"FF88C6DA", x"003B13BD", x"FFAD92AE", x"FFFAFDAA", x"00C5B837", x"001FFE23", x"FFFF169C", x"FFF505EA", x"FE7F8642", x"FDCDF990", x"FDBDF660", x"FCB63680", x"FCDC61D4", x"FBF2B188", x"FD87E390", x"FDCAB808", x"FCE2C31C", x"FC2C2E40", x"FC6C82B4", x"FC10690C", x"FD4A00EC", x"FF0DD140", x"FFC2F22F", x"00E101C7", x"FFF3FA62", x"014958D8", x"FFA217D6", x"FF8766AB", x"00C52C8B", x"FFC6B7D6", x"0053B282", x"FFCC06A9", x"FF31158D", x"FFF00A3B", x"00744C5F", x"0085CEE2", x"0059ECA2", x"FEF2B20C", x"FF3FDAD2", x"FEA96BBE", x"FE16753C", x"FE3B9E26", x"FE0AF364", x"FE503B58", x"FD6EECA8", x"FDCD2474", x"FCCD6078", x"FDAC760C", x"FFB7539A", x"FFBEBDAF", x"01E04B12", x"025A7A8C", x"01795BD8", x"00B4C118", x"00746000", x"00B26E44", x"FF20E098", x"FFB12693", x"FF4DBF4D", x"FEF75E9C", x"FF2EAA14", x"FF4358EB", x"00D5701F", x"009DFF61", x"FF29BC62", x"FF0316EF", x"011371B0", x"008410D3", x"00FD25F1", x"010F388E", x"005C7626", x"FFEDB1E5", x"006ABD2C", x"FE674706", x"FF326149", x"019EF0EE", x"020B8034", x"02F48880", x"03603EA4", x"01E71B16", x"012B0738", x"005F8B07", x"FF938EE6", x"0004C2FB", x"00F5F865", x"FFEC81A5", x"00A07455", x"FF6E7FA9", x"001D0750", x"FF24ACBD", x"FFE8B24E", x"003F37AA", x"FFB2F2DF", x"01641360", x"01096EAA", x"01CFF04E", x"0305C5DC", x"0333495C", x"02D8B2FC", x"03A00EC8", x"040A2BB8", x"01BA50A6", x"029A5514", x"0404A1D0", x"038E6D34", x"02B2BE10", x"02694E60", x"01D606CE", x"01F98120", x"016998D2", x"002A3FC6", x"FF1EDF32", x"002961B8", x"005019A5", x"FF91A3DE", x"0064E22B", x"FF887C84", x"00627E17", x"00D21C13", x"00A1D555", x"FFFE2E0C", x"0144A1FA", x"00116A2D", x"FF3C2210", x"013EABB4", x"019FBE24", x"013B8216", x"01E3B61E", x"018E87C0", x"0190C5FC", x"01669C78", x"000438A0", x"00FDBCF6", x"008A7D10", x"014EF06C", x"FFD811EB", x"0076E309", x"0089FE5D", x"FF98FEB7", x"FF8A99EC", x"FF42236D", x"00508D80", x"FF0A6A4F", x"FFC3F28C", x"001045F9", x"00537955", x"FF04D416", x"003AF092", x"FF8C201D", x"FFDC97B7", x"FF2B7688", x"FF17D79E", x"00227973", x"002B5B3C", x"00EE01BF", x"00FF8F71", x"00B16AC9", x"00552575", x"009E781E", x"0056EA7A", x"FECC5AE0", x"00C7AF0C", x"00286A18", x"FFC3FA25", x"FFAE9C2F", x"00EBD2C7", x"00CBFCF5", x"FFE4D2AC", x"FF92A1C7", x"FF62B3A2", x"00A8A9E7"
--  0.030701, 0.023824, 0.012186, -0.025738, -0.012009, 0.022801, 0.032149, -0.016884, 0.015175, -0.008363, 0.022656, -0.005366, -0.028408, -0.035449, -0.001400, 0.010526, -0.021053, 0.028099, 0.016940, 0.021537, 0.016455, -0.034446, -0.006548, 0.018551, 0.017679, -0.032495, -0.020244, 0.026032, -0.029569, 0.027068, -0.006891, 0.002620, 0.017417, 0.009610, -0.022962, 0.011451, -0.030909, -0.018365, -0.006696, -0.007851, 0.025026, -0.020334, 0.029191, 0.015782, 0.010547, 0.024698, -0.024811, -0.031045, 0.001135, 0.017518, 0.017973, 0.001470, 0.034157, 0.012689, 0.015432, -0.017310, 0.010894, -0.013369, -0.028852, -0.023244, -0.021608, -0.005400, -0.015076, 0.032317, 0.013991, -0.031048, -0.001173, 0.026918, -0.007062, -0.001500, 0.001387, -0.020182, -0.031298, -0.020586, -0.015363, 0.023458, -0.031578, 0.003381, -0.014440, -0.004028, -0.003241, -0.013881, 0.008241, 0.008441, -0.020509, 0.021944, 0.032216, -0.014831, 0.007240, -0.013385, 0.023958, -0.004254, -0.034591, 0.003532, 0.021334, -0.011789, -0.025242, -0.022226, -0.005714, 0.001681, -0.037029, -0.005603, 0.000603, 0.016743, 0.015675, -0.035163, -0.032045, -0.030735, 0.022072, -0.018192, 0.019715, -0.005318, -0.014716, 0.026874, -0.006899, -0.019311, -0.005676, -0.023721, -0.036959, -0.011663, -0.012285, -0.038346, 0.004341, -0.046138, -0.063414, -0.041555, -0.079006, -0.099334, -0.085663, -0.115829, -0.032751, -0.042507, -0.024847, -0.052292, 0.012211, -0.036484, -0.015148, -0.023666, -0.018299, 0.007611, -0.035418, -0.034963, 0.008153, 0.011540, -0.000781, -0.018736, -0.022629, -0.028337, -0.044776, -0.079477, -0.045351, -0.073414, -0.125998, -0.132398, -0.177171, -0.196766, -0.178064, -0.189284, -0.157145, -0.142351, -0.113996, -0.073422, -0.080616, -0.070510, 0.008417, -0.004146, 0.020821, 0.026859, 0.015621, -0.012211, -0.006763, -0.003048, -0.003432, -0.015386, -0.061337, -0.077592, -0.058514, -0.096431, -0.112024, -0.050237, -0.051522, -0.000374, 0.095243, 0.063766, 0.049842, 0.043894, -0.032159, -0.088303, -0.066551, -0.097592, -0.125324, -0.092968, -0.046010, -0.015672, -0.030045, -0.013794, 0.012071, -0.033499, -0.034334, 0.004749, -0.008855, -0.070672, -0.095896, -0.065840, -0.075012, -0.120191, -0.035033, 0.018048, 0.115895, 0.177350, 0.287232, 0.353330, 0.294813, 0.141802, 0.080521, 0.017030, -0.085020, -0.123095, -0.136083, -0.106383, -0.066728, -0.042212, -0.036631, 0.021979, 0.034867, 0.029158, 0.019081, 0.005002, -0.039438, -0.076573, -0.089644, -0.079761, -0.078105, -0.062137, -0.031285, 0.033375, 0.097405, 0.164169, 0.190087, 0.195717, 0.132396, 0.074693, 0.001263, -0.008069, -0.076439, -0.058722, -0.122198, -0.099994, -0.016712, -0.029304, -0.011500, 0.018041, -0.030919, -0.009397, -0.006266, -0.009582, -0.035374, -0.063461, -0.070640, -0.040871, 0.007429, 0.004031, 0.070688, 0.114255, 0.047121, 0.068631, 0.044039, -0.017257, 0.007367, 0.013595, 0.026851, 0.017509, -0.008858, -0.022497, -0.083916, -0.056733, -0.006805, -0.030808, 0.004271, -0.018714, 0.013025, 0.010166, 0.020984, -0.013080, -0.003887, 0.013481, 0.020358, 0.000318, 0.094186, 0.069153, 0.134108, 0.072005, 0.025999, -0.069602, -0.115153, -0.057441, -0.046216, 0.000248, 0.041658, 0.082787, 0.066326, 0.020805, -0.007887, -0.015174, -0.011598, 0.017897, 0.018037, -0.018864, -0.005547, 0.015254, 0.022489, -0.039143, -0.019814, 0.017828, 0.102476, 0.135709, 0.109538, 0.118234, 0.119044, 0.044654, -0.065927, -0.116933, -0.083035, -0.016155, 0.042710, 0.114683, 0.120029, 0.182560, 0.104916, 0.052733, 0.043247, -0.014837, -0.043451, 0.013454, -0.015743, 0.034418, -0.010432, -0.027712, -0.030494, -0.002502, 0.016430, 0.093338, 0.100919, 0.099075, 0.133072, 0.099443, 0.079949, -0.005546, -0.098276, -0.055838, 0.010809, 0.068547, 0.116037, 0.199886, 0.188691, 0.211887, 0.112263, 0.095085, -0.006436, -0.037146, 0.011619, 0.023873, -0.013585, 0.031240, 0.004021, 0.012494, -0.004443, -0.006881, 0.023435, 0.045886, 0.121626, 0.127033, 0.145984, 0.059860, 0.065460, -0.005858, -0.014515, 0.010985, 0.107627, 0.141675, 0.202214, 0.191646, 0.219545, 0.172492, 0.049993, 0.058302, 0.009409, -0.055188, -0.051024, -0.004383, 0.027370, 0.010261, 0.004965, -0.002479, -0.036573, 0.027374, 0.056651, 0.030708, 0.061504, 0.109227, 0.070017, 0.042160, 0.041924, 0.010702, 0.034288, 0.006527, 0.047456, 0.086991, 0.198140, 0.225913, 0.147053, 0.050164, -0.008532, -0.057123, -0.034356, -0.014566, -0.044698, -0.030645, 0.025906, 0.004793, -0.016856, 0.023116, -0.029940, -0.013602, 0.011339, 0.026960, 0.034540, 0.057589, 0.050178, 0.063542, 0.038293, 0.010770, 0.017265, -0.011010, -0.026198, 0.003601, 0.170702, 0.144802, 0.046765, -0.036152, -0.036851, -0.054678, -0.103688, -0.046676, -0.009145, 0.001219, -0.002216, -0.016961, -0.025211, -0.035233, -0.001443, -0.013039, 0.017161, -0.013927, 0.018602, -0.019558, 0.075098, 0.048810, 0.081661, 0.042148, 0.012152, -0.049288, -0.046422, 0.011761, 0.146029, 0.109353, -0.041952, -0.064469, -0.089829, -0.082625, -0.047407, -0.056425, -0.044465, -0.025203, 0.002901, -0.005341, -0.025579, 0.000960, 0.019365, -0.001559, 0.014662, -0.038543, -0.008729, -0.019549, -0.018257, 0.031710, 0.044872, -0.006014, -0.040713, -0.057373, -0.065635, 0.075252, 0.078564, 0.003054, -0.049043, -0.067501, -0.062800, -0.066081, -0.098768, -0.076046, -0.012337, 0.026980, 0.029204, 0.013964, 0.033934, -0.016411, -0.002298, -0.035465, -0.039669, -0.065512, -0.089782, -0.058527, -0.060636, -0.052188, -0.036997, -0.096123, -0.099266, -0.046945, -0.031001, 0.056314, 0.019325, -0.057206, -0.054685, -0.058221, -0.057639, -0.084393, -0.047382, -0.017707, 0.001215, -0.009885, -0.033347, 0.034928, 0.009939, 0.031505, 0.010963, -0.007516, -0.003053, -0.025509, -0.074805, -0.093172, -0.125891, -0.123627, -0.137784, -0.155855, -0.098292, -0.043631, 0.006517, -0.018610, -0.039394, -0.089921, -0.043180, -0.070337, -0.075876, -0.046314, -0.079371, -0.019462, -0.030613, -0.004216, -0.014222, 0.028872, -0.026546, 0.006409, -0.001037, -0.042832, 0.006058, -0.034856, -0.103654, -0.149536, -0.135802, -0.155121, -0.204742, -0.193097, -0.170966, -0.051968, -0.067063, -0.083570, -0.064796, -0.056096, -0.054559, -0.025693, -0.001875, -0.037046, -0.022785, -0.019142, -0.026796, 0.005797, -0.018966, 0.020667, -0.024635, -0.029239, -0.008145, 0.019297, -0.043900, -0.046947, -0.070538, -0.123121, -0.126314, -0.135441, -0.154834, -0.168180, -0.148379, -0.112844, -0.091377, -0.113847, -0.125376, -0.081352, -0.074695, -0.018371, -0.033475, -0.016680, -0.020307, 0.017771, -0.031399, -0.014554, 0.007212, -0.010062, -0.000611, 0.024136, 0.003905, -0.000111, -0.001340, -0.046933, -0.068607, -0.070561, -0.102757, -0.098098, -0.126624, -0.077162, -0.069004, -0.097319, -0.119607, -0.111754, -0.122997, -0.084716, -0.029563, -0.007453, 0.027467, -0.001468, 0.040203, -0.011463, -0.014722, 0.024069, -0.006992, 0.010217, -0.006344, -0.025258, -0.001948, 0.014197, 0.016334, 0.010977, -0.032874, -0.023455, -0.041819, -0.059759, -0.055222, -0.061163, -0.052706, -0.080209, -0.068708, -0.099930, -0.072698, -0.008871, -0.007966, 0.058630, 0.073545, 0.046064, 0.022065, 0.014206, 0.021781, -0.027237, -0.009625, -0.021759, -0.032304, -0.025554, -0.023029, 0.026054, 0.019287, -0.026155, -0.030873, 0.033624, 0.016121, 0.030902, 0.033108, 0.011287, -0.002235, 0.013030, -0.049893, -0.025100, 0.050652, 0.063904, 0.092350, 0.105499, 0.059461, 0.036502, 0.011663, -0.013238, 0.000581, 0.030026, -0.002380, 0.019587, -0.017761, 0.003544, -0.026773, -0.002845, 0.007717, -0.009406, 0.043466, 0.032401, 0.056633, 0.094455, 0.100011, 0.088953, 0.113288, 0.126242, 0.053994, 0.081339, 0.125565, 0.111136, 0.084319, 0.075355, 0.057376, 0.061707, 0.044140, 0.005157, -0.027481, 0.005051, 0.009778, -0.013472, 0.012315, -0.014589, 0.012023, 0.025648, 0.019755, -0.000222, 0.039628, 0.002126, -0.023910, 0.038900, 0.050750, 0.038514, 0.059047, 0.048649, 0.048923, 0.043776, 0.000515, 0.030974, 0.016905, 0.040886, -0.004874, 0.014513, 0.016845, -0.012574, -0.014331, -0.023176, 0.009833, -0.029979, -0.007331, 0.001986, 0.010190, -0.030661, 0.007195, -0.014145, -0.004322, -0.025944, -0.028340, 0.004208, 0.005293, 0.029054, 0.031196, 0.021657, 0.010394, 0.019344, 0.010610, -0.037554, 0.024375, 0.004933, -0.007327, -0.009935, 0.028787, 0.024901, -0.003318, -0.013351, -0.019201, 0.020589
--  Sum of weights (converted): FFFFFFFF918181A6
    );

    attribute rom_style : string;
    attribute rom_style of weights_n0 : constant is "block";
    attribute rom_style of weights_n1 : constant is "block";
    attribute rom_style of weights_n2 : constant is "block";
    attribute rom_style of weights_n3 : constant is "block";
    attribute rom_style of weights_n4 : constant is "block";
    attribute rom_style of weights_n5 : constant is "block";
    attribute rom_style of weights_n6 : constant is "block";
    attribute rom_style of weights_n7 : constant is "block";
    attribute rom_style of weights_n8 : constant is "block";
    attribute rom_style of weights_n9 : constant is "block";

begin

    read_n0 : process(clk) is
    begin
        if rising_edge(clk) then
            dout((1*DATA_WIDTH-1) downto (0*DATA_WIDTH)) <= weights_n0(to_integer(unsigned(addr)));
        end if;
    end process read_n0;

    read_n1 : process(clk) is
    begin
        if rising_edge(clk) then
            dout((2*DATA_WIDTH-1) downto (1*DATA_WIDTH)) <= weights_n1(to_integer(unsigned(addr)));
        end if;
    end process read_n1;

    read_n2 : process(clk) is
    begin
        if rising_edge(clk) then
            dout((3*DATA_WIDTH-1) downto (2*DATA_WIDTH)) <= weights_n2(to_integer(unsigned(addr)));
        end if;
    end process read_n2;

    read_n3 : process(clk) is
    begin
        if rising_edge(clk) then
            dout((4*DATA_WIDTH-1) downto (3*DATA_WIDTH)) <= weights_n3(to_integer(unsigned(addr)));
        end if;
    end process read_n3;

    read_n4 : process(clk) is
    begin
        if rising_edge(clk) then
            dout((5*DATA_WIDTH-1) downto (4*DATA_WIDTH)) <= weights_n4(to_integer(unsigned(addr)));
        end if;
    end process read_n4;

    read_n5 : process(clk) is
    begin
        if rising_edge(clk) then
            dout((6*DATA_WIDTH-1) downto (5*DATA_WIDTH)) <= weights_n5(to_integer(unsigned(addr)));
        end if;
    end process read_n5;

    read_n6 : process(clk) is
    begin
        if rising_edge(clk) then
            dout((7*DATA_WIDTH-1) downto (6*DATA_WIDTH)) <= weights_n6(to_integer(unsigned(addr)));
        end if;
    end process read_n6;

    read_n7 : process(clk) is
    begin
        if rising_edge(clk) then
            dout((8*DATA_WIDTH-1) downto (7*DATA_WIDTH)) <= weights_n7(to_integer(unsigned(addr)));
        end if;
    end process read_n7;

    read_n8 : process(clk) is
    begin
        if rising_edge(clk) then
            dout((9*DATA_WIDTH-1) downto (8*DATA_WIDTH)) <= weights_n8(to_integer(unsigned(addr)));
        end if;
    end process read_n8;

    read_n9 : process(clk) is
    begin
        if rising_edge(clk) then
            dout((10*DATA_WIDTH-1) downto (9*DATA_WIDTH)) <= weights_n9(to_integer(unsigned(addr)));
        end if;
    end process read_n9;

end rtl;