-- VHDL Memory Module for Layer Weights: test_weights
-- Number of Neurons: 10
-- Number of Inputs per Neuron: 784
-- Data Width: 32 bits
-- Address Width: 10 bits
-- Expected Data Encoding: fixed_point
-- Res for 0x02000000 : ['0000000040000000', '000000005E000000', '0000000068000000', 'FFFFFFFFB8000000', 'FFFFFFFFC0000000', '0000000068000000', 'FFFFFFFF9C000000', '0000000034000000', 'FFFFFFFF98000000', '000000004C000000']
-- Res from input file mnist_sample_input.npz with label [2]: 0x['0000000009441262', 'FFFFFFFFBE133CFE', '000000004E3896F2', '0000000062DB7DFF', 'FFFFFFFFF2C7B377', 'FFFFFFFFA893E5C6', 'FFFFFFFFAF45DF4E', '0000000020AC5BA9', '00000000040D5587', '0000000008DB120C']
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity test_weights is
    port(
        clk   : in  std_logic;
        addr  : in  std_logic_vector(9 downto 0); -- Same addr for all neurons within a layer
        dout  : out std_logic_vector(32*10-1 downto 0) -- DATA_WIDTH * N_NEURONS -> 320 bits
    );
end test_weights;

architecture rtl of test_weights is
    constant DATA_WIDTH : integer := 32;
    constant N_INPUTS  : integer := 784;
   type weight_array is array (0 to N_INPUTS-1) of std_logic_vector(DATA_WIDTH-1 downto 0);
    constant weights_n0 : weight_array := (
     x"8030C6A9", x"80C534EE", x"011DD0E0", x"803AAF12", x"007434D5", x"81053D94", x"00A86C6E", x"805AED2B", x"80DE8CFA", x"002AC7D9", x"008DBD5C", x"00FD30C3", x"80B2BA2C", x"80907B76", x"0037C086", x"004F57AE", x"00707C50", x"00A095D0", x"80425777", x"00A28B37", x"00D7B5E1", x"804C6D0B", x"00D026EE", x"008EF1C5", x"0102103E", x"80A642BE", x"80907973", x"80549802", x"000ED750", x"00AF99E1", x"80A704A3", x"00927A20", x"8068DBC2", x"00B0B9FE", x"800E1822", x"8101007E", x"80A23E43", x"80D5D706", x"008EE4CF", x"80C46CDC", x"8016F0C8", x"003D6CEE", x"80A520AA", x"0052D06D", x"811BF1FE", x"80D1769B", x"810B068A", x"805A27BD", x"806C23E2", x"0029429B", x"80364532", x"008985B4", x"010C3A68", x"0068F8D7", x"8073437E", x"8111F5AE", x"0069F84E", x"8090F4F3", x"0094E1B9", x"00C41585", x"0070D56F", x"01125680", x"01141CE0", x"003B811A", x"80DC561D", x"00F433D9", x"80A420AC", x"80A96607", x"00CAF9DC", x"00AA3BBE", x"000C8050", x"80429DB7", x"814AED9A", x"807205B7", x"00CAC040", x"00098E01", x"8011B12F", x"805414C8", x"8072883B", x"00A9690E", x"00109FC2", x"00BE0A32", x"8033C8E4", x"007FD3C0", x"0078C3C2", x"002EA797", x"00B7D756", x"00B87C7A", x"010E995A", x"00DAA9F4", x"8057B59C", x"810FC3A4", x"00102B73", x"804C560A", x"80B0A146", x"809BE93A", x"807C98E4", x"002DB3DB", x"8073D081", x"814CE7BC", x"81715464", x"815E5632", x"81949D52", x"00069DBC", x"8027C763", x"00803C77", x"8050C2CE", x"0016C22E", x"00589B7B", x"8116F10E", x"0019DAC1", x"801391F2", x"80A40807", x"80E30550", x"0102F954", x"00EE907B", x"0083D2B3", x"00FFBF02", x"80A95998", x"80832FA2", x"800F661C", x"80E0EEB3", x"810E865A", x"81B81E1E", x"804238FA", x"80C0D9D8", x"00418587", x"019673EC", x"8034F1DB", x"8071295B", x"00502D7C", x"80F5459D", x"80BB6C3F", x"0065863A", x"80FD945D", x"81283DB6", x"80D40FCD", x"805E5537", x"808D6445", x"8097E002", x"00762EC0", x"0031B80B", x"805DD134", x"80E37E60", x"806C2FBB", x"80B6457A", x"80CDD767", x"81C08AB4", x"80CD5BE2", x"82078710", x"81DDE10E", x"8168FDBA", x"00A275A5", x"009DBAB5", x"01988E0C", x"035D9988", x"03198088", x"02DE3AAC", x"0080DF37", x"000635C4", x"8051543A", x"009A9B3E", x"807F4A96", x"8192031E", x"807A2CD3", x"81118A86", x"804B19A5", x"80514C85", x"00FD4493", x"005A9E00", x"8033E7A1", x"002A2170", x"80789CCE", x"001E79BA", x"80342985", x"80BD9020", x"81CAF0D2", x"805C6B93", x"80ED87F8", x"8078E835", x"015A6748", x"027E0CD0", x"03464844", x"03099DBC", x"02EF7C5C", x"044A86B8", x"0431E240", x"01160E0A", x"011AF556", x"8012020D", x"002F7EF5", x"80441514", x"811D0D22", x"808C4476", x"0063DA0A", x"8033D6E3", x"80F5B212", x"00E9D38C", x"8096E0CB", x"802E79F6", x"80250FB3", x"8092D514", x"81F3D410", x"80AC7FA0", x"81DB2882", x"817BD8BA", x"8011AD39", x"8057696B", x"0056A738", x"00FBE8BA", x"017476B8", x"02089EC4", x"03104790", x"0489ACA0", x"034CEDA0", x"0252C940", x"01AD8FA6", x"013B6298", x"01467F9A", x"810AC07C", x"80A105E6", x"800D4D9C", x"0073AF1B", x"810FF4BC", x"806E58D7", x"80FC3F64", x"80C30924", x"007EF2D4", x"80967FED", x"803B6C10", x"81A2A12E", x"80F21788", x"81A56698", x"80165260", x"80A73A41", x"00203677", x"0008A8E0", x"0162A602", x"02D6D3C0", x"02B9E4EC", x"026E8458", x"03B22818", x"03ED5738", x"024FFFF4", x"02F772DC", x"0161B1E0", x"01A24138", x"003E6F18", x"81310130", x"80911378", x"003FB3CB", x"003F2527", x"808D3DDB", x"011A9FA8", x"803A0C56", x"80E67CB2", x"810C18C8", x"005B795C", x"80CE1678", x"80DED000", x"8121B404", x"80A25C8A", x"80CFC99E", x"80360A20", x"02204334", x"02B2AE28", x"0277AB10", x"0020ACC4", x"01D896C6", x"0148E324", x"03CFCB60", x"042290F8", x"0356D18C", x"02E9F288", x"03279488", x"01E378FA", x"009905F4", x"810047EE", x"005C5C88", x"805FF839", x"8005598D", x"81013692", x"805ACFF2", x"80D6F28E", x"80EBDDC0", x"81609D3A", x"816EC26A", x"801724CE", x"007F286E", x"0105A0C6", x"010A6732", x"00D7F568", x"0093C33D", x"0177CC2C", x"007B6ADB", x"825F7B00", x"815166D8", x"00933A4C", x"01C73F2E", x"022832D4", x"04193330", x"03B99054", x"04AE6F78", x"02727CE0", x"017F0EC8", x"812446D4", x"0104B2A6", x"807CDDA8", x"00AFFE32", x"0038C6EA", x"003BE520", x"806A6D83", x"801FC7F9", x"80E6BA4D", x"80C24FB1", x"00315D76", x"0125D776", x"800D9E41", x"016F7DE4", x"0166E378", x"01D0F0BA", x"8006A1A3", x"828D5E78", x"85254710", x"85D7CFD0", x"834A34B8", x"815944E6", x"02B965B8", x"021CACA8", x"04A9E008", x"0619BF78", x"04BE7B38", x"01D9EAAC", x"813C7E64", x"010C5D36", x"80325DF8", x"81117510", x"011FAF40", x"8083AC16", x"804E4E2B", x"007EC8DC", x"80B27B9E", x"00592060", x"017FBA04", x"009122A0", x"016C7C4A", x"013A61CA", x"01C8056E", x"809C29A4", x"83A45EA4", x"86EC8B28", x"86C6D0C8", x"876306B8", x"86C79998", x"81CDEFDE", x"00A71CC3", x"02A91E84", x"03970F4C", x"05AE05D0", x"05C1EF38", x"02B1BBF0", x"80E1F249", x"0105C004", x"00167F5B", x"008CB750", x"00E39A78", x"00F2A6E5", x"811599C8", x"009A6126", x"000AA447", x"0211A434", x"0168B39E", x"0190397A", x"0259B650", x"02A08C04", x"00BE9101", x"82107268", x"849D5960", x"87407EF0", x"88530BE0", x"88735E90", x"861B85E0", x"83CB65A0", x"8096B484", x"01D72226", x"03068C08", x"0470C770", x"04C7DF88", x"01A03A74", x"000DB3F5", x"8045C7D1", x"002CE58F", x"00BE4C4B", x"80616395", x"00E58711", x"00B59BC8", x"8124EAD8", x"00BA82F6", x"02033D9C", x"02A54958", x"0297828C", x"034B2F98", x"0262D1FC", x"80F82749", x"8496B140", x"87E04D08", x"8802A7D0", x"8A0E9A70", x"89F478A0", x"860D1690", x"836AB080", x"00443225", x"02309350", x"047A40B0", x"03BEF2E4", x"04EA7990", x"0304553C", x"807BE62E", x"010A129C", x"00DB3E1F", x"00032E15", x"008CCD33", x"806990B1", x"8139000C", x"0038DC9B", x"02A0B8D0", x"02C7BD58", x"0488CD90", x"031E3084", x"05151B88", x"03627FDC", x"817E7708", x"86612BE8", x"87F0D9C0", x"897FB2C0", x"8957EC20", x"87E36200", x"8466F950", x"827C2844", x"80008559", x"01F079A8", x"02D259A8", x"048EA2F0", x"02E27114", x"01AE4C40", x"003EEB2E", x"805219B3", x"00C6DCA7", x"001FF70A", x"810E961E", x"80253EB7", x"80CD79AD", x"002848C7", x"02778168", x"02D8184C", x"042CE798", x"048FD2A8", x"03CAE598", x"02D73478", x"82AFC6D8", x"85850108", x"882719C0", x"8A18F710", x"88473310", x"85855F48", x"83E655F0", x"81224902", x"022DA33C", x"0289F73C", x"019B2754", x"037EF2B0", x"026655B8", x"0000FE33", x"000BE2CF", x"0056557A", x"8058A36B", x"0065C7E0", x"80FA4DDC", x"00C291FA", x"009C9546", x"00AE6279", x"02B03AA0", x"0453D9B0", x"03A62ED8", x"0475E130", x"041CB6C0", x"01358BA4", x"83194B5C", x"84B05330", x"869A2D90", x"88D62620", x"861271B8", x"834F30B4", x"0016B394", x"01428F32", x"024F946C", x"00FB1B05", x"02720F38", x"0315ACBC", x"0078C4B8", x"8056D516", x"002A3325", x"009A4006", x"808F4842", x"00203372", x"8000912D", x"00405825", x"811E993A", x"00853FCD", x"02C8C570", x"029B530C", x"04460C10", x"04AB3BB0", x"0499CEC0", x"035089B8", x"80D2E701", x"843F6958", x"8471BCE0", x"85C192F8", x"83E46E30", x"814FD6B0", x"808151F9", x"0110CE8C", x"003D1770", x"00EC2183", x"013A6920", x"0169C118", x"803F8DAF", x"80F82C16", x"007464DF", x"00F6DA5F", x"8104AB56", x"006C5DE0", x"80D68A5A", x"00043303", x"008C6A73", x"00A6CF5C", x"00A0BA7A", x"03643138", x"04183ED8", x"0427DC60", x"057BC980", x"02A72DC4", x"006DFD3A", x"81EDDAAE", x"8262802C", x"81EF4BEA", x"80F72DFF", x"804FFFEC", x"007729FC", x"012116BC", x"809C877B", x"0026C33B", x"00A0622E", x"000F4029", x"00775757", x"8011473C", x"00B70592", x"801D4FAE", x"80B8FECC", x"00CEB785", x"002B954B", x"805F2C0C", x"8132DD4C", x"00112B5D", x"80190B20", x"0225E62C", x"02FEF18C", x"0260095C", x"0391FC8C", x"0339C858", x"03707208", x"01BB1A92", x"801E0BCE", x"00F2B16C", x"00589B72", x"8015EC08", x"0110E580", x"00659ECC", x"00D87348", x"800DD5CD", x"01067FDA", x"008C3510", x"007FB7C7", x"815650C2", x"00E00B72", x"80FBEC6E", x"010649B6", x"800C1FE8", x"81036BD6", x"00468A94", x"808961A2", x"813F4FFC", x"0024E1DC", x"01596F1E", x"02A32B14", x"021EC5B0", x"04632FB0", x"046F4320", x"03D90748", x"02B9F154", x"00EE35FB", x"00B1D1F5", x"013346D0", x"000120A0", x"807568BE", x"806AFAD6", x"815B2CC4", x"80ED0839", x"80B63F47", x"80A5D93E", x"80F9AC66", x"801377FA", x"8030A928", x"00552A41", x"000D3A85", x"80921A03", x"8064BC11", x"8008C550", x"80E05023", x"8043D26D", x"001245FC", x"0154DB8E", x"01AF802E", x"030C0680", x"032D9C5C", x"034A6618", x"0527A5C8", x"03A52F78", x"03E05C64", x"02BF88E4", x"01A5B59C", x"006398E6", x"00C2588F", x"8048AC8B", x"80A112EF", x"001C17DA", x"81D593AA", x"804C3AE8", x"0085B6E6", x"00B1E04A", x"80EBDE0C", x"006854CE", x"80A6A5EF", x"800B6E90", x"803D0D0B", x"80F5A6D3", x"8125DB20", x"80F5F8FF", x"0056F2B8", x"0097FBEB", x"807244A3", x"00A594FB", x"01EF2BA2", x"01D7D1F4", x"04368888", x"04C0F758", x"03509B98", x"0138FB10", x"0115A74A", x"000517E0", x"8031B293", x"81F581B8", x"82487E08", x"8086C893", x"80931C55", x"80B0A2CC", x"8099E0A6", x"809DE713", x"00EC284A", x"8032B55D", x"00D3012C", x"010529EE", x"00250FD2", x"003D9D16", x"8016D2E9", x"00B94DEA", x"812F1B38", x"0031DA06", x"80A99E6B", x"800CFB86", x"80B29C8A", x"8119BC8A", x"80C66926", x"002BB963", x"813D398C", x"8172E3A8", x"8155C0B8", x"81CD984A", x"80F7A8E5", x"8072B2FA", x"81074674", x"00705201", x"80E17063", x"80D68E6F", x"8095FA32", x"80CCFB27", x"80CC5E18", x"8104B14E", x"81034CCC", x"004C5C59", x"00B26D05", x"0112A4CA", x"00F8CC44", x"80150635", x"0025B1EA", x"80DE850E", x"001183C7", x"81BA8282", x"8060F7AA", x"81039212", x"80F7956B", x"80F8A962", x"81D64AEC", x"80483391", x"80A33F30", x"805D1884", x"80D14321", x"0003E0B6", x"0054057A", x"00369DCE", x"00ADCCB3", x"804C9E8E", x"00B72456", x"0040F051", x"00B00615", x"011CF638", x"00423FC0", x"806C97C5", x"801D1C17", x"00525E00", x"00314D52", x"8050BD8B", x"00DE1B00", x"009DF52A", x"80D4847E", x"804D2BE8", x"806D942B", x"811B3ECC", x"80423800", x"80C2F3E8", x"8105FD24", x"80D1E0AF", x"80D69E28", x"00B20531", x"00173287", x"00DC51C3", x"0029806C", x"0027557C", x"0065EBC4", x"00286AB8", x"80E7A317", x"80AD1425", x"8046ED91", x"000465F6", x"006E3745", x"0070A775", x"00E819D1", x"003B8F40", x"8063DA47", x"80DC0C20", x"80D713DD", x"80B08EC6", x"0055FC49", x"009A98F4", x"00FA31D2", x"806264F1", x"801DF87E", x"8064B5C7", x"80145584", x"004218D5", x"801E02F6", x"8007D581", x"0010CB5E", x"005D747F", x"8060B982", x"80B357F9", x"004171EF", x"8029955D", x"8085E91C", x"007ADE82", x"0002A742", x"802A8F0D", x"808DA10C"
--  -0.005954, -0.024073, 0.034890, -0.007164, 0.014185, -0.031890, 0.020560, -0.011099, -0.027167, 0.005222, 0.017302, 0.030907, -0.021817, -0.017637, 0.006806, 0.009685, 0.013731, 0.019603, -0.008098, 0.019842, 0.026332, -0.009329, 0.025409, 0.017449, 0.031502, -0.020295, -0.017636, -0.010326, 0.001812, 0.021436, -0.020388, 0.017880, -0.012800, 0.021573, -0.001720, -0.031372, -0.019805, -0.026104, 0.017443, -0.023978, -0.002800, 0.007498, -0.020157, 0.010109, -0.034661, -0.025569, -0.032596, -0.011005, -0.013201, 0.005037, -0.006625, 0.016787, 0.032743, 0.012814, -0.014070, -0.033442, 0.012936, -0.017695, 0.018174, 0.023936, 0.013774, 0.033489, 0.033705, 0.007264, -0.026897, 0.029810, -0.020035, -0.020679, 0.024777, 0.020780, 0.001526, -0.008132, -0.040397, -0.013919, 0.024750, 0.001166, -0.002160, -0.010264, -0.013981, 0.020680, 0.002029, 0.023198, -0.006321, 0.015604, 0.014742, 0.005695, 0.022442, 0.022520, 0.033032, 0.026692, -0.010707, -0.033174, 0.001974, -0.009318, -0.021561, -0.019032, -0.015210, 0.005579, -0.014138, -0.040638, -0.045084, -0.042766, -0.049391, 0.000808, -0.004856, 0.015654, -0.009859, 0.002778, 0.010816, -0.034050, 0.003156, -0.002389, -0.020023, -0.027712, 0.031613, 0.029122, 0.016092, 0.031219, -0.020673, -0.016014, -0.001880, -0.027458, -0.033023, -0.053725, -0.008084, -0.023541, 0.007998, 0.049616, -0.006463, -0.013814, 0.009787, -0.029940, -0.022879, 0.012393, -0.030955, -0.036162, -0.025886, -0.011515, -0.017260, -0.018539, 0.014427, 0.006069, -0.011452, -0.027770, -0.013206, -0.022250, -0.025127, -0.054754, -0.025068, -0.063419, -0.058335, -0.044066, 0.019831, 0.019254, 0.049872, 0.105176, 0.096863, 0.089628, 0.015731, 0.000758, -0.009928, 0.018873, -0.015538, -0.049074, -0.014914, -0.033391, -0.009168, -0.009924, 0.030916, 0.011062, -0.006336, 0.005143, -0.014723, 0.003720, -0.006367, -0.023140, -0.056023, -0.011282, -0.028995, -0.014759, 0.042286, 0.077887, 0.102329, 0.094924, 0.091734, 0.134097, 0.131089, 0.033942, 0.034541, -0.002198, 0.005798, -0.008311, -0.034796, -0.017122, 0.012189, -0.006328, -0.029992, 0.028543, -0.018418, -0.005673, -0.004524, -0.017924, -0.061014, -0.021057, -0.058003, -0.046368, -0.002158, -0.010670, 0.010578, 0.030751, 0.045467, 0.063552, 0.095737, 0.141806, 0.103141, 0.072606, 0.052437, 0.038499, 0.039856, -0.032562, -0.019656, -0.001624, 0.014122, -0.033198, -0.013470, -0.030792, -0.023808, 0.015497, -0.018372, -0.007254, -0.051102, -0.029552, -0.051441, -0.002725, -0.020414, 0.003932, 0.001057, 0.043292, 0.088724, 0.085192, 0.075991, 0.115498, 0.122722, 0.072266, 0.092706, 0.043176, 0.051056, 0.007621, -0.037232, -0.017709, 0.007776, 0.007708, -0.017241, 0.034500, -0.007086, -0.028136, -0.032727, 0.011166, -0.025157, -0.027199, -0.035364, -0.019820, -0.025365, -0.006597, 0.066438, 0.084312, 0.077108, 0.003989, 0.057689, 0.040147, 0.119116, 0.129220, 0.104348, 0.091058, 0.098582, 0.059018, 0.018680, -0.031284, 0.011275, -0.011715, -0.000653, -0.031398, -0.011085, -0.026239, -0.028792, -0.043044, -0.044770, -0.002825, 0.015522, 0.031937, 0.032520, 0.026362, 0.018037, 0.045874, 0.015066, -0.074155, -0.041187, 0.017972, 0.055572, 0.067407, 0.128076, 0.116402, 0.146293, 0.076476, 0.046760, -0.035678, 0.031823, -0.015242, 0.021484, 0.006931, 0.007311, -0.012992, -0.003880, -0.028165, -0.023720, 0.006026, 0.035869, -0.001662, 0.044860, 0.043810, 0.056755, -0.000809, -0.079757, -0.160800, -0.182594, -0.102808, -0.042147, 0.085132, 0.066000, 0.145737, 0.190643, 0.148252, 0.057851, -0.038634, 0.032759, -0.006148, -0.033381, 0.035118, -0.016073, -0.009559, 0.015477, -0.021787, 0.010880, 0.046842, 0.017717, 0.044493, 0.038377, 0.055667, -0.019063, -0.113815, -0.216375, -0.211769, -0.230838, -0.211865, -0.056389, 0.020399, 0.083144, 0.112190, 0.177493, 0.179924, 0.084196, -0.027581, 0.031952, 0.002746, 0.017177, 0.027784, 0.029621, -0.033887, 0.018845, 0.001299, 0.064653, 0.044031, 0.048856, 0.073451, 0.082098, 0.023263, -0.064508, -0.144208, -0.226623, -0.260137, -0.264083, -0.190860, -0.118579, -0.018397, 0.057511, 0.094549, 0.138767, 0.149399, 0.050809, 0.001673, -0.008518, 0.005481, 0.023230, -0.011888, 0.028019, 0.022169, -0.035757, 0.022768, 0.062896, 0.082677, 0.080995, 0.102928, 0.074563, -0.030292, -0.143395, -0.246130, -0.250324, -0.314283, -0.311093, -0.189098, -0.106774, 0.008325, 0.068430, 0.139923, 0.117059, 0.153622, 0.094279, -0.015124, 0.032480, 0.026763, 0.000388, 0.017188, -0.012886, -0.038208, 0.006941, 0.082119, 0.086882, 0.141700, 0.097435, 0.158827, 0.105774, -0.046688, -0.199362, -0.248151, -0.296838, -0.291983, -0.246507, -0.137570, -0.077656, -0.000064, 0.060605, 0.088178, 0.142412, 0.090142, 0.052527, 0.007681, -0.010022, 0.024275, 0.003902, -0.033031, -0.004547, -0.025082, 0.004918, 0.077088, 0.088879, 0.130482, 0.142557, 0.118518, 0.088770, -0.083957, -0.172486, -0.254773, -0.315547, -0.258691, -0.172531, -0.121867, -0.035435, 0.068071, 0.079342, 0.050190, 0.109247, 0.074992, 0.000121, 0.001451, 0.010539, -0.010820, 0.012424, -0.030555, 0.023751, 0.019114, 0.021287, 0.084012, 0.135236, 0.114036, 0.139390, 0.128505, 0.037786, -0.096838, -0.146524, -0.206321, -0.276141, -0.189751, -0.103417, 0.002771, 0.039375, 0.072214, 0.030653, 0.076423, 0.096396, 0.014742, -0.010600, 0.005151, 0.018829, -0.017491, 0.003931, -0.000069, 0.007855, -0.034985, 0.016266, 0.087008, 0.081460, 0.133551, 0.145902, 0.143775, 0.103581, -0.025745, -0.132741, -0.138884, -0.179880, -0.121635, -0.040996, -0.015786, 0.033302, 0.007457, 0.028825, 0.038380, 0.044159, -0.007758, -0.030294, 0.014208, 0.030133, -0.031820, 0.013228, -0.026189, 0.000513, 0.017141, 0.020363, 0.019620, 0.105981, 0.127960, 0.129866, 0.171361, 0.082908, 0.013426, -0.060285, -0.074524, -0.060461, -0.030173, -0.009766, 0.014546, 0.035289, -0.019108, 0.004732, 0.019578, 0.001862, 0.014568, -0.002109, 0.022342, -0.003578, -0.022582, 0.025234, 0.005320, -0.011618, -0.037459, 0.002096, -0.003057, 0.067126, 0.093621, 0.074223, 0.111571, 0.100804, 0.107476, 0.054090, -0.003668, 0.029626, 0.010816, -0.002676, 0.033313, 0.012405, 0.026422, -0.001689, 0.032043, 0.017115, 0.015591, -0.041787, 0.027349, -0.030752, 0.032018, -0.001480, -0.031668, 0.008611, -0.016770, -0.038979, 0.004502, 0.042167, 0.082418, 0.066256, 0.137108, 0.138582, 0.120243, 0.085198, 0.029078, 0.021707, 0.037509, 0.000138, -0.014332, -0.013059, -0.042380, -0.028935, -0.022247, -0.020245, -0.030478, -0.002377, -0.005940, 0.010396, 0.001615, -0.017835, -0.012297, -0.001071, -0.027382, -0.008279, 0.002231, 0.041609, 0.052673, 0.095218, 0.099318, 0.102832, 0.161090, 0.113914, 0.121138, 0.085881, 0.051478, 0.012158, 0.023724, -0.008871, -0.019662, 0.003429, -0.057321, -0.009305, 0.016323, 0.021713, -0.028792, 0.012736, -0.020343, -0.001395, -0.007453, -0.029987, -0.035871, -0.030026, 0.010614, 0.018553, -0.013949, 0.020213, 0.060446, 0.057595, 0.131657, 0.148555, 0.103590, 0.038206, 0.033893, 0.000622, -0.006067, -0.061219, -0.071349, -0.016453, -0.017958, -0.021562, -0.018784, -0.019275, 0.028828, -0.006190, 0.025757, 0.031880, 0.004524, 0.007521, -0.002786, 0.022620, -0.037000, 0.006085, -0.020705, -0.001585, -0.021803, -0.034392, -0.024220, 0.005337, -0.038724, -0.045275, -0.041718, -0.056347, -0.030232, -0.014001, -0.032138, 0.013711, -0.027519, -0.026191, -0.018308, -0.025022, -0.024947, -0.031823, -0.031653, 0.009321, 0.021781, 0.033526, 0.030371, -0.002566, 0.004601, -0.027163, 0.002138, -0.054017, -0.011837, -0.031686, -0.030223, -0.030354, -0.057409, -0.008814, -0.019928, -0.011364, -0.025545, 0.000473, 0.010257, 0.006667, 0.021216, -0.009353, 0.022356, 0.007927, 0.021487, 0.034785, 0.008087, -0.013256, -0.003553, 0.010055, 0.006018, -0.009856, 0.027112, 0.019282, -0.025942, -0.009420, -0.013376, -0.034576, -0.008083, -0.023798, -0.031981, -0.025620, -0.026198, 0.021731, 0.002832, 0.026894, 0.005066, 0.004802, 0.012442, 0.004934, -0.028276, -0.021128, -0.008658, 0.000537, 0.013454, 0.013752, 0.028333, 0.007270, -0.012189, -0.026861, -0.026255, -0.021552, 0.010496, 0.018872, 0.030541, -0.012011, -0.003659, -0.012294, -0.002482, 0.008068, -0.003664, -0.000956, 0.002050, 0.011408, -0.011807, -0.021893, 0.007989, -0.005076, -0.016347, 0.014999, 0.000324, -0.005195, -0.017289
--  Sum of weights (converted): 000000005AF884A0
    );

    constant weights_n1 : weight_array := (
     x"80267E10", x"80F8C7E5", x"00428EA2", x"000463F9", x"00B18B03", x"0012E436", x"00176449", x"004FB345", x"00DEA0EC", x"808A41C3", x"00AEAAAA", x"00478D3E", x"80C33595", x"00656D51", x"80AFE25B", x"805C1D04", x"808B75AE", x"80C70A5E", x"00E66BC1", x"810581A8", x"00924A45", x"8107515A", x"80239B92", x"00117319", x"00CFFDFC", x"8069E135", x"005435C9", x"002D5230", x"00AC2505", x"001164D2", x"006D8D42", x"80B0BD5E", x"80CB5033", x"0104B290", x"80D53F3E", x"803214C3", x"80257CC6", x"011BD0CE", x"80410109", x"80E0D1EA", x"804C4D47", x"00944590", x"0075B2A9", x"00F68FED", x"803FF42D", x"0086480F", x"8115183C", x"00703AFE", x"0085A5D5", x"00BC47D1", x"80A7E5FE", x"804E1EED", x"0046C820", x"80CFE7D3", x"80E8BC2A", x"8119775C", x"00105509", x"00B5AEEE", x"004B265C", x"0011CF8B", x"0065C3F8", x"80B7EA70", x"001E6484", x"804AE897", x"80986FF0", x"00EECB2C", x"80F5F456", x"0015B8FB", x"8113AE7C", x"801042C8", x"8081A100", x"006F3DE8", x"80AB0CE2", x"009DA854", x"8111D6A2", x"008FA8FA", x"80F6798D", x"008B40B9", x"80853CBA", x"80049642", x"8036D43F", x"00BDA1BC", x"005FE23B", x"8101D0B4", x"001AE630", x"80C9D583", x"00DACCF0", x"00300349", x"804B617C", x"8096C89A", x"00607910", x"80BFDE13", x"005F1491", x"00526BAD", x"003CA6E7", x"804B6483", x"8199883A", x"0055D94A", x"80C86205", x"80B51C14", x"80A70F14", x"00164A34", x"001B38DC", x"807D3C1E", x"000EDADA", x"8158EB30", x"80226CDF", x"8115A992", x"0058259C", x"80D2C684", x"8069478E", x"00CC843E", x"01179BFC", x"80AFA7C5", x"80A21937", x"002427E4", x"007289EC", x"803440EC", x"80730991", x"8106B060", x"8007FD1A", x"004F8968", x"816C7DB4", x"8005B26B", x"00DBA772", x"020E2CD4", x"011CB224", x"00EC9880", x"010F4C84", x"00A78034", x"01682E1A", x"00E3F228", x"020F3878", x"022849C4", x"800E0E5F", x"006F2AFD", x"8052EC6C", x"00AD0370", x"808631A9", x"0013C8C2", x"00AF0C73", x"810C0798", x"80F69215", x"8094231F", x"00BA08B8", x"00AF8969", x"8111671E", x"8070FFC8", x"81CEADB6", x"82324F40", x"80B4B446", x"807B4569", x"0006CAED", x"01D46B66", x"01C6DF64", x"011146DC", x"80B325EE", x"81271462", x"01399220", x"02013300", x"0329DE98", x"01E68E8C", x"01C62604", x"012A20B4", x"009B567E", x"002566E6", x"0117D4DC", x"800189C9", x"003E49A0", x"0115F9FC", x"011B126A", x"807A9796", x"00FA9AAF", x"002E23DF", x"80B9DD45", x"8034FFFD", x"829CA4AC", x"8216A460", x"81E99392", x"832315CC", x"81BA0890", x"81008DD0", x"8038F104", x"826EDB78", x"82E21050", x"81DD0190", x"006C834E", x"01E4D464", x"02882550", x"01AADEB4", x"8075F1B5", x"812FBECC", x"80636619", x"00C92161", x"0001B234", x"801C7A40", x"80C69447", x"8091674B", x"80E279A3", x"00E338BD", x"804AFB9D", x"817054EC", x"80E2AF5B", x"819FD160", x"82E77B88", x"8346A978", x"83963C9C", x"84FBE758", x"834B39A8", x"8102D8F0", x"81E8B10A", x"82F78DAC", x"81CA8D94", x"825C46EC", x"81577BB8", x"8002FDF2", x"80AAD131", x"005DF340", x"81432B5C", x"81D22428", x"81DCD5A2", x"002AC704", x"803FAC1F", x"8021F1FC", x"804C41A1", x"808D7844", x"0031C3B0", x"00D65169", x"80D04643", x"807E142B", x"820E8F00", x"828673F0", x"820559EC", x"840DBF28", x"83B5345C", x"84CB6EF0", x"839E8E58", x"81744322", x"01970AEA", x"8039E391", x"80005F9D", x"805EB4CA", x"803C317B", x"805524C7", x"8205D008", x"819768D8", x"8332F5C4", x"82553944", x"80834AB6", x"804B5971", x"803F68E8", x"8045B0EF", x"80B2D626", x"00B1CBA1", x"800D04D4", x"8016CB67", x"001BBDB7", x"00480D1D", x"81B8A93C", x"823A95BC", x"8210A2BC", x"832D21C0", x"851E5AB0", x"85AC5890", x"82BAEDC4", x"010062BE", x"03DB7BE4", x"05653A88", x"016B4E12", x"00B92C3C", x"81CEC4BA", x"81B36CEE", x"82499574", x"82CEEF88", x"81B198F6", x"82A8924C", x"8236FFD8", x"8199248C", x"00A72679", x"0064C917", x"80D67C57", x"008DFD74", x"0107A24C", x"812D5EC0", x"00AEDFC2", x"804F1B59", x"80EC3224", x"809B3295", x"8173B450", x"830655EC", x"8367C9B4", x"8429C3F0", x"82CE529C", x"00890037", x"07610120", x"07818E68", x"043AB960", x"00084810", x"8217A224", x"83F19700", x"842A34E8", x"81F79C02", x"81690BC2", x"80B1CF2A", x"8116EF4C", x"80754FA5", x"80567E06", x"00C88CB5", x"807E5FC8", x"00B815B9", x"00C79BD8", x"8114A850", x"8017B0F8", x"8093DD93", x"817A0B54", x"80F83BB1", x"827B9440", x"828AFDA8", x"8558BC60", x"84DDDE48", x"84B0EEF8", x"020B2B18", x"0A8A3B00", x"0B8D9BC0", x"0428EBC8", x"82361950", x"82B6D258", x"840B1E40", x"82C19F5C", x"82CD2A18", x"817CCE96", x"001A8A55", x"816604B8", x"8134DFF0", x"002E950A", x"00285020", x"8035859C", x"00FF4F3C", x"80B1C5E4", x"80B6D5FC", x"80EC151B", x"808BF446", x"81029226", x"809DF2A1", x"82593F48", x"834BFF50", x"85CEB820", x"85899AB0", x"839990B4", x"02E26678", x"0CC07750", x"099FB670", x"024E1100", x"83A00104", x"84443080", x"8224913C", x"83399FE0", x"80710B2A", x"80B644DF", x"0073AA1C", x"80CF1969", x"00B012B7", x"001EF254", x"001669D3", x"00C7C0F5", x"81162A98", x"80EC8E6D", x"01180C80", x"80BE3D40", x"81261574", x"80CA0361", x"81C70B9A", x"828493A0", x"84C7E828", x"85A73730", x"88485D20", x"84C3F7B0", x"06A07A50", x"0DAC64B0", x"091B06A0", x"804F4CF6", x"84D827A0", x"84BAAF40", x"83924EC8", x"82ACE8CC", x"81CB1392", x"005480F2", x"80B5CCBC", x"001BC212", x"00B50870", x"801CA7B9", x"809E1E68", x"80C63B00", x"806BD815", x"0068268C", x"80F6567F", x"80310E31", x"0014E200", x"0018B789", x"812F79EA", x"824980E0", x"8372A1A8", x"85BB8520", x"86D87878", x"838ED10C", x"07154330", x"0C3EA7A0", x"069DA518", x"8321D84C", x"86466000", x"846A4D50", x"82840470", x"828F6A14", x"826DB4CC", x"8182703C", x"812503E2", x"0054EF2B", x"80D6AF29", x"801FE356", x"803E1BD4", x"80B19286", x"0084990E", x"8078F242", x"80112BB9", x"80E2C0D2", x"8090BE89", x"80DBD3C5", x"81B9BD06", x"830E5E28", x"83D6CB60", x"860D0608", x"85C7A278", x"80E35ECE", x"08E41D50", x"0A850970", x"04D57498", x"85AE87B0", x"871D2DF8", x"84E94638", x"833D5BDC", x"827BBB3C", x"80CA4BC7", x"81C10DBE", x"804700AF", x"80611C21", x"810F30C4", x"80793C46", x"0049B16D", x"0037E3B9", x"00D4BB2A", x"00C4F1D5", x"80A80FED", x"80A371E1", x"80DC7ACC", x"822EBF48", x"8260BBA8", x"83CFD184", x"837BA524", x"83531FB4", x"8240A670", x"016B7FDE", x"08859EE0", x"0976AF90", x"01777FFE", x"859D1848", x"864E5B50", x"840461E0", x"8310C24C", x"823809CC", x"81DF026A", x"809B2A08", x"805960DE", x"817919F8", x"80E2DB08", x"80013D3C", x"006E40EE", x"008E563C", x"80ADD176", x"81247E6E", x"801C9908", x"805EC450", x"809A8901", x"8236EA80", x"81AF483E", x"82EF4A08", x"8248FEE8", x"82A4E6AC", x"0099DD22", x"043959A8", x"081A7D80", x"07A1BEF8", x"8151FFA4", x"842A9700", x"85D37560", x"84BED880", x"82E7F7FC", x"824C8634", x"8135C75C", x"807B857B", x"81BFCE44", x"00381B24", x"806D9551", x"80507F49", x"0039FE32", x"00E4C6FE", x"809F0FB9", x"80C8E642", x"009FF650", x"80E78E98", x"80E5A184", x"82A01958", x"82A8792C", x"81E3D132", x"826A516C", x"80CEEE04", x"02512388", x"047C2DF8", x"062EED90", x"0367A180", x"00595643", x"8445D1B0", x"8528A358", x"84B1FAC0", x"834EC7B0", x"81A7F5CC", x"81B43C6E", x"804BDFBB", x"80F8B63F", x"80AF64EC", x"0076EFF3", x"800DB493", x"80399DF3", x"0061CF63", x"00E69E16", x"00430AE4", x"00ADF4CD", x"0049533D", x"811F179E", x"82175DB4", x"82779F94", x"820C39D0", x"003E4188", x"01A8D232", x"025A8964", x"0292ECB8", x"04708E88", x"0156C46E", x"005882C1", x"8259A744", x"831905AC", x"8365E388", x"835B5148", x"8124FA9C", x"820103E4", x"80D15D9C", x"800FBBE8", x"816C9718", x"80087627", x"806B6517", x"00D03447", x"80BA47DA", x"00B16353", x"00AF2069", x"007D06DF", x"00AAA233", x"80F5DDA7", x"82B41100", x"80EBED45", x"80D6C7BE", x"0041C04E", x"801912D7", x"00B19B79", x"803D3F8A", x"019A70CA", x"017B8E3C", x"006CCE28", x"80EC3864", x"831AE174", x"82DB9290", x"82856028", x"822902B8", x"806900B2", x"808CD9D8", x"005B6FBC", x"805806EB", x"81189574", x"80576C6D", x"00CDB735", x"00B229EA", x"005A86E8", x"805C7F72", x"8125ECFC", x"80CCEDF8", x"0065BE5D", x"809EA673", x"00824AB5", x"00D91E58", x"006C8A2A", x"01310FD8", x"815EA848", x"8220E56C", x"8213EDBC", x"814C98B2", x"0078DA37", x"0000FEC4", x"81A17CA6", x"80CB37D0", x"8292E5F4", x"825EE068", x"81A70F42", x"81288BF8", x"8094B263", x"80677B60", x"007DB893", x"8102ED90", x"002B1497", x"00051C20", x"004D495A", x"011E8DAA", x"00A73783", x"809C1308", x"8047014D", x"00C916C4", x"00DE82CC", x"020E12E0", x"013F181A", x"008998D1", x"821ECF4C", x"83D583E8", x"827A3BA4", x"002BD592", x"012BEF82", x"020B08F4", x"80846839", x"000C48AE", x"819EC8F2", x"81C9AFA0", x"80E61580", x"0008F787", x"008AD94E", x"0031F0E7", x"8019E25E", x"800FD19E", x"80769A5E", x"801A412D", x"80143704", x"00F82B94", x"00A1081D", x"80D4F4F0", x"00B25A0E", x"00AEB4FC", x"019709AC", x"00DC0227", x"01586478", x"8191E0C4", x"816D85D0", x"81F96FDA", x"828D310C", x"80F27AF4", x"01B29DA8", x"01499F30", x"011D722A", x"8109235A", x"0004BE69", x"8163A27E", x"80F3B0F4", x"80D4534B", x"006AB79C", x"80117051", x"81190EF8", x"80A6048D", x"80876533", x"810F74DA", x"0025767D", x"006831AD", x"803AF5E3", x"807BD8A2", x"0024D149", x"80A99030", x"80B84B78", x"808D4355", x"802BB3FB", x"82949030", x"826294C4", x"836EC080", x"82D3467C", x"82D455F0", x"801F296F", x"00539311", x"807D3B6F", x"005C7F34", x"00B185EE", x"0061DEBF", x"007D394B", x"8129A726", x"811D119E", x"80E39526", x"005C7BCF", x"80FCDD64", x"80DF5535", x"808DCF6A", x"810DA8A8", x"00006448", x"00298266", x"80B22BBA", x"00AB4598", x"809EC2C8", x"80C592FA", x"0021500D", x"802014D7", x"81AF34FE", x"827AA3A8", x"822BB8FC", x"81742C8C", x"80BAF388", x"8098905B", x"813FE1CA", x"817C6DC6", x"81348DC6", x"807C8601", x"800E0F4E", x"808CA4C1", x"80EC669D", x"001C8D01", x"80E90976", x"80E0AE75", x"80EDD9E7", x"804F4772", x"01026A86", x"00725F30", x"8022B09D", x"003C198D", x"007274B0", x"8002F401", x"80F77C4D", x"80CC21CB", x"80ED67B8", x"803D3BFF", x"8156E926", x"808C93B3", x"80C99594", x"00B1CA5B", x"009340EB", x"006DAE1F", x"801947D7", x"80786DC2", x"003C1028", x"80D2A593", x"8081B95A", x"803D8E6A", x"8045BF62", x"81157A7A", x"00744673", x"00F0E50A", x"80A15FE7", x"004EDE0E", x"8021EE47", x"800AABB9", x"00110DD2", x"00FD898C", x"00272DB5", x"80B95A46", x"8069DFB8", x"008E2EF1", x"005A2954", x"0003F410", x"802A6B3F", x"8074BCB7", x"806C3641", x"809F6E04", x"002ACEE5", x"004DDDC8", x"00DBBFAF", x"80464826", x"0011E72D", x"00BC568E", x"007EB9F0", x"002568B9", x"0059A793", x"000F2BD9", x"80FAF723", x"000B4769", x"803FF330", x"0108051A"
--  -0.004699, -0.030369, 0.008125, 0.000536, 0.021673, 0.002306, 0.002855, 0.009729, 0.027176, -0.016877, 0.021322, 0.008734, -0.023829, 0.012381, -0.021470, -0.011244, -0.017024, -0.024297, 0.028128, -0.031922, 0.017858, -0.032143, -0.004347, 0.002130, 0.025390, -0.012925, 0.010280, 0.005532, 0.021014, 0.002123, 0.013373, -0.021575, -0.024819, 0.031823, -0.026031, -0.006113, -0.004576, 0.034645, -0.007935, -0.027444, -0.009314, 0.018100, 0.014367, 0.030098, -0.007807, 0.016392, -0.033825, 0.013700, 0.016314, 0.022983, -0.020495, -0.009536, 0.008640, -0.025379, -0.028410, -0.034359, 0.001994, 0.022178, 0.009174, 0.002174, 0.012423, -0.022451, 0.003710, -0.009144, -0.018608, 0.029150, -0.030024, 0.002652, -0.033653, -0.001985, -0.015824, 0.013579, -0.020880, 0.019245, -0.033428, 0.017537, -0.030087, 0.016999, -0.016264, -0.000560, -0.006693, 0.023148, 0.011705, -0.031472, 0.003284, -0.024638, 0.026709, 0.005861, -0.009202, -0.018406, 0.011776, -0.023421, 0.011606, 0.010061, 0.007404, -0.009203, -0.049992, 0.010480, -0.024461, -0.022108, -0.020393, 0.002721, 0.003323, -0.015287, 0.001813, -0.042104, -0.004202, -0.033894, 0.010760, -0.025729, -0.012852, 0.024965, 0.034132, -0.021442, -0.019787, 0.004414, 0.013982, -0.006379, -0.014043, -0.032067, -0.000975, 0.009709, -0.044494, -0.000695, 0.026813, 0.064230, 0.034753, 0.028881, 0.033118, 0.020447, 0.043967, 0.027825, 0.064358, 0.067418, -0.001716, 0.013570, -0.010123, 0.021120, -0.016381, 0.002415, 0.021368, -0.032718, -0.030099, -0.018083, 0.022709, 0.021428, -0.033374, -0.013794, -0.056479, -0.068641, -0.022059, -0.015048, 0.000829, 0.057180, 0.055526, 0.033359, -0.021869, -0.036020, 0.038278, 0.062646, 0.098861, 0.059394, 0.055438, 0.036393, 0.018962, 0.004566, 0.034159, -0.000188, 0.007603, 0.033933, 0.034555, -0.014965, 0.030591, 0.005632, -0.022689, -0.006470, -0.081621, -0.065264, -0.059763, -0.098033, -0.053959, -0.031318, -0.006951, -0.076032, -0.090096, -0.058228, 0.013246, 0.059183, 0.079119, 0.052108, -0.014397, -0.037078, -0.012134, 0.024552, 0.000207, -0.003476, -0.024241, -0.017749, -0.027646, 0.027737, -0.009153, -0.044962, -0.027672, -0.050759, -0.090757, -0.102376, -0.112089, -0.155750, -0.102933, -0.031598, -0.059655, -0.092719, -0.055976, -0.073764, -0.041929, -0.000365, -0.020852, 0.011469, -0.039449, -0.056902, -0.058207, 0.005222, -0.007773, -0.004144, -0.009309, -0.017269, 0.006075, 0.026162, -0.025424, -0.015390, -0.064277, -0.078913, -0.063153, -0.126678, -0.115870, -0.149833, -0.113105, -0.045442, 0.049688, -0.007067, -0.000046, -0.011561, -0.007348, -0.010394, -0.063210, -0.049733, -0.099971, -0.072903, -0.016027, -0.009198, -0.007740, -0.008507, -0.021831, 0.021704, -0.001589, -0.002783, 0.003386, 0.008795, -0.053792, -0.069651, -0.064531, -0.099259, -0.159955, -0.177288, -0.085318, 0.031297, 0.120542, 0.168607, 0.044349, 0.022604, -0.056490, -0.053153, -0.071482, -0.087761, -0.052929, -0.083078, -0.069214, -0.049944, 0.020404, 0.012303, -0.026182, 0.017333, 0.032182, -0.036788, 0.021347, -0.009657, -0.028833, -0.018945, -0.045374, -0.094523, -0.106419, -0.130098, -0.087686, 0.016724, 0.230591, 0.234565, 0.132168, 0.001011, -0.065385, -0.123241, -0.130152, -0.061476, -0.044073, -0.021705, -0.034050, -0.014320, -0.010558, 0.024481, -0.015427, 0.022471, 0.024366, -0.033772, -0.002892, -0.018050, -0.046148, -0.030302, -0.077585, -0.079467, -0.167082, -0.152084, -0.146598, 0.063863, 0.329374, 0.361036, 0.129995, -0.069104, -0.084817, -0.126357, -0.086136, -0.087544, -0.046485, 0.003240, -0.043703, -0.037704, 0.005686, 0.004921, -0.006533, 0.031166, -0.021701, -0.022319, -0.028819, -0.017084, -0.031564, -0.019281, -0.073394, -0.103027, -0.181484, -0.173047, -0.112496, 0.090137, 0.398494, 0.300746, 0.072030, -0.113282, -0.133324, -0.066964, -0.100784, -0.013799, -0.022250, 0.014119, -0.025281, 0.021493, 0.003778, 0.002736, 0.024384, -0.033956, -0.028877, 0.034186, -0.023223, -0.035899, -0.024660, -0.055548, -0.078684, -0.149403, -0.176662, -0.258833, -0.148922, 0.207090, 0.427294, 0.284549, -0.009680, -0.151386, -0.147789, -0.111610, -0.083607, -0.056040, 0.010315, -0.022192, 0.003388, 0.022099, -0.003498, -0.019302, -0.024198, -0.013165, 0.012714, -0.030071, -0.005988, 0.002549, 0.003017, -0.037045, -0.071473, -0.107743, -0.179141, -0.213925, -0.111184, 0.221346, 0.382648, 0.206744, -0.097881, -0.196091, -0.137976, -0.078615, -0.080007, -0.075892, -0.047173, -0.035768, 0.010368, -0.026207, -0.003893, -0.007582, -0.021676, 0.016186, -0.014764, -0.002096, -0.027680, -0.017669, -0.026834, -0.053923, -0.095504, -0.119970, -0.189090, -0.180619, -0.027755, 0.277846, 0.328740, 0.151057, -0.177555, -0.222312, -0.153476, -0.101240, -0.077604, -0.024694, -0.054816, -0.008667, -0.011854, -0.033104, -0.014799, 0.008996, 0.006822, 0.025968, 0.024041, -0.020515, -0.019952, -0.026914, -0.068206, -0.074308, -0.119118, -0.108843, -0.103897, -0.070392, 0.044372, 0.266311, 0.295738, 0.045837, -0.175427, -0.197065, -0.125535, -0.095796, -0.069341, -0.058473, -0.018941, -0.010910, -0.046033, -0.027692, -0.000151, 0.013459, 0.017375, -0.021218, -0.035705, -0.003491, -0.011568, -0.018864, -0.069204, -0.052647, -0.091710, -0.071411, -0.082630, 0.018782, 0.132001, 0.253234, 0.238494, -0.041260, -0.130199, -0.182063, -0.148297, -0.090816, -0.071841, -0.037815, -0.015078, -0.054664, 0.006849, -0.013377, -0.009826, 0.007079, 0.027927, -0.019417, -0.024524, 0.019527, -0.028266, -0.028031, -0.082043, -0.083066, -0.059060, -0.075478, -0.025260, 0.072405, 0.140159, 0.193229, 0.106400, 0.010905, -0.133523, -0.161211, -0.146726, -0.103367, -0.051753, -0.053251, -0.009262, -0.030360, -0.021410, 0.014519, -0.001673, -0.007033, 0.011940, 0.028152, 0.008184, 0.021235, 0.008951, -0.035045, -0.065352, -0.077102, -0.063992, 0.007600, 0.051858, 0.073552, 0.080435, 0.138740, 0.041842, 0.010805, -0.073444, -0.096804, -0.106188, -0.104897, -0.035764, -0.062624, -0.025557, -0.001921, -0.044506, -0.001033, -0.013110, 0.025416, -0.022739, 0.021654, 0.021378, 0.015262, 0.020829, -0.030013, -0.084481, -0.028800, -0.026218, 0.008026, -0.003061, 0.021681, -0.007477, 0.050103, 0.046332, 0.013282, -0.028835, -0.097031, -0.089303, -0.078781, -0.067506, -0.012818, -0.017194, 0.011162, -0.010745, -0.034251, -0.010672, 0.025112, 0.021749, 0.011051, -0.011291, -0.035880, -0.025016, 0.012420, -0.019366, 0.015905, 0.026504, 0.013249, 0.037239, -0.042805, -0.066516, -0.064933, -0.040600, 0.014752, 0.000121, -0.050963, -0.024807, -0.080432, -0.074082, -0.051643, -0.036200, -0.018151, -0.012632, 0.015347, -0.031607, 0.005259, 0.000624, 0.009434, 0.034980, 0.020412, -0.019052, -0.008668, 0.024547, 0.027162, 0.064218, 0.038952, 0.016797, -0.066261, -0.119814, -0.077421, 0.005351, 0.036613, 0.063847, -0.016163, 0.001500, -0.050633, -0.055870, -0.028086, 0.001095, 0.016949, 0.006096, -0.003160, -0.001931, -0.014478, -0.003205, -0.002468, 0.030294, 0.019657, -0.025996, 0.021771, 0.021327, 0.049687, 0.026856, 0.042040, -0.049057, -0.044619, -0.061699, -0.079735, -0.029600, 0.053054, 0.040237, 0.034844, -0.032365, 0.000579, -0.043412, -0.029747, -0.025919, 0.013027, -0.002129, -0.034309, -0.020266, -0.016528, -0.033137, 0.004573, 0.012719, -0.007197, -0.015118, 0.004494, -0.020699, -0.022497, -0.017244, -0.005335, -0.080635, -0.074534, -0.107270, -0.088290, -0.088420, -0.003804, 0.010202, -0.015287, 0.011291, 0.021670, 0.011947, 0.015286, -0.036335, -0.034798, -0.027781, 0.011290, -0.030867, -0.027262, -0.017311, -0.032917, 0.000048, 0.005067, -0.021749, 0.020907, -0.019380, -0.024118, 0.004066, -0.003916, -0.052638, -0.077471, -0.067837, -0.045431, -0.022821, -0.018624, -0.039048, -0.046439, -0.037665, -0.015201, -0.001716, -0.017168, -0.028858, 0.003485, -0.028447, -0.027427, -0.029035, -0.009678, 0.031545, 0.013961, -0.004235, 0.007336, 0.013972, -0.000360, -0.030211, -0.024918, -0.028980, -0.007475, -0.041859, -0.017160, -0.024607, 0.021703, 0.017975, 0.013389, -0.003086, -0.014701, 0.007332, -0.025714, -0.015835, -0.007514, -0.008514, -0.033872, 0.014194, 0.029406, -0.019699, 0.009627, -0.004142, -0.001303, 0.002082, 0.030949, 0.004783, -0.022626, -0.012924, 0.017356, 0.011006, 0.000483, -0.005178, -0.014250, -0.013209, -0.019462, 0.005226, 0.009505, 0.026825, -0.008579, 0.002185, 0.022990, 0.015470, 0.004567, 0.010944, 0.001852, -0.030635, 0.001377, -0.007806, 0.032229
--  Sum of weights (converted): FFFFFFFE96129AAF
    );

    constant weights_n2 : weight_array := (
     x"01081546", x"003A0B1E", x"01058054", x"8096AE0A", x"00FE4B9E", x"00FBE651", x"800B2EB0", x"80EACA95", x"805E6967", x"804E3DD9", x"0004D52B", x"810942A0", x"00363ECC", x"8075CDE3", x"8046A8AF", x"8096EF0A", x"803DC592", x"810FB7EC", x"809B1CAC", x"001AF400", x"00BFB70C", x"0109DFA8", x"80DD513A", x"007ADB60", x"80A4EBDA", x"80E23423", x"800CE22B", x"80A7D527", x"80FBF9E1", x"81116B2E", x"80C3D50C", x"00F06A9A", x"00A3256F", x"8073E245", x"80C48E4A", x"80E351A3", x"80AE4D38", x"807D411D", x"00A7835D", x"00544DDF", x"807C5510", x"00C60159", x"80B223EE", x"80EC05BD", x"004E7D4A", x"80A19796", x"004D7C6C", x"00F2B83B", x"808E446C", x"80CE7453", x"006D597A", x"810863F2", x"01050696", x"808A2B2E", x"008D7250", x"80E8A501", x"80C60845", x"00203A64", x"0067FAD0", x"00E2C9D9", x"00F3D44A", x"8010F469", x"8027B439", x"002AD87D", x"804A66FB", x"000303F1", x"812703B4", x"81018C34", x"00B8B3C2", x"80C54CFA", x"00D0C246", x"00117CE5", x"002FBFF5", x"00D41E76", x"80EFF95D", x"8082FA40", x"800A0A2B", x"0035C9C5", x"813B15F8", x"005D660C", x"80AB4859", x"00291582", x"00C5F06A", x"801D2502", x"80094164", x"8015DC0D", x"00F42729", x"00A60B38", x"00302408", x"80A9AF59", x"808E9227", x"0122602E", x"014B9D72", x"019C266C", x"00779CBC", x"02948120", x"01CD3158", x"02DDB8C4", x"02BEFC20", x"019515D0", x"00AAD806", x"01955D9C", x"80C29FEE", x"0032EA15", x"81B571B4", x"80DED3F4", x"815B5220", x"80B6B8F7", x"006AB659", x"80D25E28", x"80FD8564", x"00D132EC", x"009C2E3E", x"800339AE", x"80CE69A7", x"804DD51E", x"805E6C6B", x"00DE29AE", x"00166FF4", x"00A5C076", x"00ED8A55", x"02558C44", x"0462E188", x"0558C580", x"0560FB08", x"04D41780", x"06563C98", x"04FC5270", x"03BEC7B0", x"02605180", x"00F1F536", x"00476020", x"8084021C", x"805092DC", x"80F9E7B6", x"005B8F4C", x"80BABF31", x"80934C7E", x"806DE007", x"8112DF20", x"80C00E3C", x"8108BD94", x"80115155", x"00038B78", x"8043B089", x"80688FD6", x"021BE848", x"01B69E18", x"03C0BB58", x"0534EBD0", x"0472C700", x"05731B48", x"06566DC0", x"06E38DA8", x"05C61698", x"06B64190", x"0483FDA8", x"0347ED1C", x"02E89CD4", x"00081398", x"0038AD53", x"81240B44", x"81A2AD6E", x"000F447C", x"0078C096", x"8006D23C", x"80B6AAA2", x"800D3515", x"808CB3DA", x"00D52E73", x"000D17AF", x"003EDF3C", x"00C922DB", x"00ED2EEE", x"00DD2296", x"03AB3C78", x"042FCFC8", x"033BD558", x"04CA41F8", x"03FDD70C", x"0346ACB4", x"02A1EBEC", x"03494C94", x"024AD518", x"03B99E90", x"031B52D4", x"00C8E79F", x"01084018", x"8140E388", x"80FCEA16", x"82114DC8", x"8171E872", x"804DDA9A", x"003DAC2A", x"8013F435", x"809498EA", x"00CC80BC", x"00C0D16B", x"0033D102", x"8086605B", x"0066AD19", x"00BD0499", x"02EF1C20", x"028EBCE4", x"0290218C", x"022BDE04", x"02997C58", x"02004C94", x"02A30E44", x"0232F72C", x"00B32373", x"0124DA7E", x"80129E51", x"8097098C", x"000DFE7C", x"8034237D", x"80DDC971", x"0045D48E", x"819CF7EE", x"82198FF8", x"813AE580", x"805DCB2D", x"8027CE01", x"01064BAA", x"807BA37A", x"80982B9A", x"001A54E5", x"00D61EC4", x"0078DD26", x"01731B36", x"01BE9748", x"02577BEC", x"018DE1C0", x"016F3A20", x"00FDC8F6", x"00214C84", x"00065D99", x"00BF396B", x"017ED23C", x"0052C37F", x"0179FDE2", x"00941779", x"800ECBA0", x"8030E053", x"80CE9CBA", x"004A4226", x"810DC6C8", x"80E04619", x"823158E8", x"810ECB6E", x"00103B59", x"00E8F5CD", x"008B1E90", x"0036C8A9", x"8121DDEC", x"0005A55C", x"808D4BC5", x"803EB317", x"00B8490C", x"8124A6AE", x"805F807C", x"81B42640", x"803030BD", x"803AB2F2", x"82701938", x"8119F788", x"81088B8A", x"00CAB6F0", x"01FC3064", x"008A5769", x"0007BF9E", x"00C8F8E4", x"80561FC0", x"80E6C628", x"803B091D", x"8216D6E8", x"812D0326", x"0061BBA5", x"0063BEB5", x"80BE617E", x"004BC626", x"80E03D05", x"80A0B955", x"00BF3424", x"805546B7", x"809836E4", x"80B4ED68", x"8238BC68", x"84013408", x"84071208", x"847E78C8", x"83C8EF10", x"858FB860", x"84C56730", x"836DB750", x"81F995D8", x"80017054", x"8023A93D", x"80301734", x"800C2864", x"814BC6F8", x"81B342B2", x"80567644", x"81403CCC", x"8147DAD0", x"804A403B", x"00D01211", x"80F4F9FB", x"809B3BF9", x"80D485F9", x"80196141", x"80199C36", x"8124248E", x"8039164C", x"839B370C", x"837E9DDC", x"863510F0", x"85D9F2F8", x"86236688", x"87BCDF88", x"86BFBCE0", x"880887B0", x"855CC650", x"836FF66C", x"808968B6", x"003D04B4", x"009D7DD6", x"00433E30", x"80E5BE2B", x"00294DDC", x"817C030E", x"80B22FB2", x"812D0F8E", x"80982736", x"80F5E1EC", x"010D0E2A", x"00307FED", x"80D29600", x"0016B06A", x"809EEBDC", x"806CDC4D", x"818B9628", x"84B18890", x"85A9D958", x"87228128", x"86A58A08", x"88AD5980", x"87FB9740", x"86E9DF28", x"861D2DA0", x"851EB8C8", x"82A16C54", x"814B2DA0", x"81A167A6", x"80743298", x"0042249A", x"008E4D12", x"805A92D0", x"8293BC98", x"81EC7242", x"812E383A", x"0086CC2B", x"8105F8FE", x"00693D74", x"80504E04", x"0069A694", x"0059EEA7", x"80B0CF09", x"8016AC0F", x"81F9C99C", x"85698840", x"848162E8", x"84C48BA8", x"85280250", x"86154A48", x"8516C7E8", x"856481E8", x"849F3CD8", x"83170CD0", x"82C0B6C0", x"8233B74C", x"82EF3F7C", x"800E062C", x"80FE1875", x"8007015F", x"80DAB034", x"81CF639E", x"80B3C81A", x"0014B620", x"00EF73DC", x"80304047", x"011C8CD0", x"004CAC45", x"00AB3F6A", x"8043FA55", x"00B78E87", x"0070BC18", x"83142BC8", x"8278A7AC", x"84636380", x"83F3972C", x"83B5B840", x"81CFA266", x"81F55BEA", x"80E856DF", x"80FEBDDC", x"80C2EEB7", x"82E816A0", x"81EBCD08", x"815E8668", x"80B305C7", x"81987CE8", x"80FCB9BB", x"82B6E368", x"830C85B8", x"81B51598", x"8109FFB8", x"01212C88", x"807BB678", x"8016641E", x"00798473", x"81029230", x"00DE9746", x"8081E121", x"80674416", x"8184B1D4", x"81AA5780", x"8159EEE2", x"813BFA36", x"00991ACF", x"00FCD4A4", x"030F5AD4", x"0357CFEC", x"0358D4FC", x"0127B98A", x"00B28433", x"01542C54", x"009D26DE", x"81857DB6", x"81214E70", x"82675300", x"815CC588", x"81CCB2FE", x"0034B259", x"0082C475", x"00E32E58", x"806646DF", x"80DBEF8C", x"002E0E23", x"8092D4E3", x"808EB51C", x"0100921E", x"00116D82", x"00576D0C", x"0217F1E4", x"01B4CE22", x"00D779C8", x"028A4FC4", x"0385A1F0", x"02EFF15C", x"04E06028", x"04025CB8", x"0209A004", x"02F0E1CC", x"0161B3C2", x"01E2B5D4", x"8052571C", x"81070376", x"00A7A64F", x"803E0F07", x"0078ABD1", x"017F13A0", x"008C2445", x"00A4FBAF", x"00F1AEBA", x"010C7B00", x"801EF56D", x"00CD0F56", x"005ED87E", x"00C7151A", x"00D6C0E0", x"039B752C", x"03827AF4", x"02EF8A10", x"0377BFC4", x"02136B34", x"03DEC6C4", x"042F5E30", x"0507A9F0", x"04946018", x"0385FBA0", x"03432E60", x"01D6AD0E", x"01115216", x"011A723C", x"00BA3889", x"00679FD6", x"02EE6E50", x"0276DBC4", x"01E63EAA", x"036E0B58", x"02802784", x"801DC607", x"009A2CC7", x"80B58390", x"0064F688", x"01005C5E", x"014A8FFE", x"02B11CB4", x"0362F410", x"044C6170", x"046A5500", x"03C7B874", x"038A57CC", x"04B1C850", x"049A1838", x"04C85650", x"03B0AD0C", x"02A0BD08", x"021234D0", x"039FE0C8", x"0230C050", x"009B2E09", x"01280574", x"0295FCE8", x"02C8A228", x"03809DCC", x"03EB0DB0", x"03724970", x"01E31652", x"004EC4CB", x"00C3FED3", x"00BB3807", x"00F00AC0", x"80231C70", x"80129C58", x"022FC184", x"02F01204", x"04ED13B8", x"047CACE8", x"04164038", x"03A9E834", x"0528F288", x"054BD570", x"053AD350", x"030D09DC", x"02A95C34", x"01D8DB64", x"00CE1ED9", x"00E2D2E2", x"02646CD4", x"01A071C4", x"03F25874", x"048B6630", x"051B8EE0", x"054589E8", x"03BF12E8", x"01E88574", x"00D5492B", x"80782306", x"809B252C", x"80368E3B", x"0091A68D", x"013BA1F6", x"02DAB938", x"02E4E9DC", x"0410BF28", x"03C952D4", x"05544678", x"03CEC5D8", x"034CA710", x"0407FD08", x"022F693C", x"00AA231D", x"802D9B6F", x"80660742", x"019933E2", x"0043BD1D", x"036E6600", x"04663190", x"043AB4E0", x"04BDC048", x"05A5C760", x"046D3010", x"03922AF0", x"01BE6FAE", x"809CD098", x"00B48373", x"00938AF9", x"80CFFC26", x"0083B98B", x"8044FF00", x"00946117", x"023D1AB8", x"02DC06FC", x"0331C2FC", x"02E880CC", x"045782A8", x"03D71C9C", x"017BD202", x"8026E4BD", x"806A2203", x"820622CC", x"81F50A7A", x"806F6BFC", x"020BD034", x"01DEF34C", x"0395E3EC", x"03597A50", x"032701BC", x"0397F060", x"02E69A60", x"016D9604", x"014CD36A", x"0085AAB6", x"00B626C6", x"00729675", x"001EAF9F", x"009946AE", x"808FD157", x"013FE0C4", x"018C17F4", x"00E66C9E", x"01B5B3EA", x"010FF352", x"00CF688F", x"01191844", x"007402F7", x"810467C0", x"8192F892", x"83696540", x"82F068D0", x"8061FB1F", x"80E1B1A6", x"01EE25F0", x"0345AE8C", x"038EDF58", x"031EF724", x"01584396", x"01B27D86", x"004E4756", x"80262D23", x"00E05B6E", x"80636E92", x"80D187F7", x"80EADBB5", x"00B641B3", x"0006DBB5", x"011D4966", x"00285D6A", x"81611E40", x"807E33A3", x"80484626", x"810EFDEE", x"81C14430", x"834AFB4C", x"83C5E484", x"82FBCB98", x"848B3988", x"832D2E34", x"82A7A6AC", x"811CA120", x"803F7F6E", x"8073A20A", x"0040C0BF", x"01EA8092", x"00E67910", x"0106081E", x"80644E88", x"00FA217B", x"803EDB6E", x"80629D80", x"003B5974", x"8068D50E", x"80768BF2", x"803C653D", x"803CBF1D", x"810ECAF8", x"8076EF5D", x"8287C038", x"8159E14C", x"81850BB2", x"82ACD2DC", x"831E6D88", x"83CFD9C0", x"8230C398", x"818F6860", x"814FF874", x"81D1D9F8", x"8110E44A", x"001330F0", x"809CA783", x"8108C10E", x"814848FA", x"00708933", x"00726CD0", x"011CBDA2", x"8085CC51", x"007FABDE", x"8060CC6B", x"8048B6D9", x"00AAB625", x"810C41AA", x"00D34C0A", x"00766C96", x"80DA3870", x"003BC905", x"80EFD5EE", x"80DA2920", x"8160FF76", x"82334F8C", x"812E839E", x"8077912F", x"811A9C1A", x"816E9984", x"80B919C5", x"808398B1", x"80F606F1", x"817469F2", x"811AD8E6", x"8085AE79", x"002BC2D3", x"00DD6728", x"800DFCB4", x"006435E8", x"00AA1617", x"807D6F82", x"80611485", x"00C2107A", x"00D17A4A", x"004553D0", x"80E22C65", x"00A3E1DC", x"80F75A25", x"0083B07B", x"0006F63E", x"00399612", x"814556EC", x"809A4C49", x"0040EFA7", x"00A5F5D3", x"808DC332", x"00D0A4D8", x"80702A0D", x"80DE5ABA", x"80A6E7D3", x"800D941B", x"804D1047", x"007AAFB6", x"80ABF101", x"80564397", x"81227100", x"00EEBBE5", x"80371D95", x"80E6A33A", x"800E1E26", x"800088B6", x"0051415E", x"80201CE9", x"00B80BC1", x"8064F62B", x"8057D41A", x"804633B9", x"003368E6", x"00E96E74", x"800EE3FE", x"00DECF60", x"00E36D10", x"809BBD58", x"801D34C5", x"808F30D8", x"007519FD", x"806B7B4F", x"0054A788", x"000ED959", x"80C10E2F", x"80C5E898", x"811E4188", x"80A462A4", x"0051AFCC", x"0011D33D", x"00DC0B28", x"81014326", x"80088CA9"
--  0.032237, 0.007085, 0.031922, -0.018394, 0.031042, 0.030749, -0.001365, -0.028661, -0.011525, -0.009551, 0.000590, -0.032380, 0.006622, -0.014380, -0.008625, -0.018425, -0.007540, -0.033169, -0.018935, 0.003290, 0.023403, 0.032455, -0.027016, 0.014997, -0.020132, -0.027613, -0.001573, -0.020487, -0.030759, -0.033376, -0.023905, 0.029348, 0.019915, -0.014146, -0.023994, -0.027749, -0.021277, -0.015290, 0.020448, 0.010291, -0.015177, 0.024171, -0.021746, -0.028811, 0.009581, -0.019726, 0.009459, 0.029629, -0.017367, -0.025202, 0.013348, -0.032274, 0.031863, -0.016866, 0.017266, -0.028399, -0.024174, 0.003934, 0.012693, 0.027684, 0.029764, -0.002070, -0.004847, 0.005230, -0.009082, 0.000368, -0.036013, -0.031439, 0.022547, -0.024085, 0.025483, 0.002135, 0.005829, 0.025893, -0.029294, -0.015988, -0.001226, 0.006566, -0.038463, 0.011401, -0.020909, 0.005015, 0.024162, -0.003558, -0.001130, -0.002668, 0.029804, 0.020269, 0.005877, -0.020713, -0.017404, 0.035446, 0.040480, 0.050311, 0.014601, 0.080628, 0.056298, 0.089566, 0.085814, 0.049449, 0.020855, 0.049483, -0.023758, 0.006215, -0.053399, -0.027201, -0.042398, -0.022305, 0.013026, -0.025680, -0.030947, 0.025537, 0.019065, -0.000394, -0.025197, -0.009501, -0.011526, 0.027119, 0.002739, 0.020233, 0.028997, 0.072943, 0.137070, 0.167086, 0.168088, 0.150890, 0.198027, 0.155801, 0.117039, 0.074258, 0.029536, 0.008713, -0.016114, -0.009836, -0.030506, 0.011177, -0.022796, -0.017981, -0.013412, -0.033554, -0.023444, -0.032317, -0.002114, 0.000433, -0.008263, -0.012764, 0.065907, 0.053542, 0.117277, 0.162710, 0.139011, 0.170301, 0.198050, 0.215278, 0.180431, 0.209748, 0.141112, 0.102530, 0.090895, 0.000986, 0.006919, -0.035650, -0.051108, 0.001864, 0.014740, -0.000833, -0.022298, -0.001612, -0.017176, 0.026023, 0.001598, 0.007675, 0.024553, 0.028953, 0.026994, 0.114653, 0.130836, 0.101054, 0.149690, 0.124736, 0.102377, 0.082266, 0.102698, 0.071635, 0.116409, 0.097085, 0.024525, 0.032257, -0.039171, -0.030873, -0.064612, -0.045155, -0.009504, 0.007528, -0.002436, -0.018139, 0.024964, 0.023537, 0.006325, -0.016403, 0.012534, 0.023073, 0.091688, 0.079924, 0.080094, 0.067855, 0.081236, 0.062537, 0.082404, 0.068721, 0.021867, 0.035749, -0.002273, -0.018437, 0.001708, -0.006365, -0.027074, 0.008524, -0.050411, -0.065620, -0.038440, -0.011449, -0.004859, 0.032019, -0.015093, -0.018575, 0.003214, 0.026138, 0.014754, 0.045301, 0.054515, 0.073179, 0.048570, 0.044828, 0.030980, 0.004065, 0.000777, 0.023343, 0.046731, 0.010103, 0.046142, 0.018078, -0.001806, -0.005966, -0.025221, 0.009065, -0.032932, -0.027377, -0.068524, -0.033056, 0.001981, 0.028438, 0.016982, 0.006687, -0.035384, 0.000689, -0.017248, -0.007654, 0.022496, -0.035724, -0.011658, -0.053241, -0.005883, -0.007165, -0.076184, -0.034420, -0.032293, 0.024745, 0.062035, 0.016887, 0.000946, 0.024533, -0.010513, -0.028171, -0.007206, -0.065288, -0.036745, 0.011930, 0.012176, -0.023240, 0.009250, -0.027373, -0.019620, 0.023340, -0.010410, -0.018581, -0.022086, -0.069426, -0.125147, -0.125863, -0.140438, -0.118278, -0.173794, -0.149097, -0.107143, -0.061717, -0.000176, -0.004353, -0.005870, -0.001484, -0.040500, -0.053132, -0.010554, -0.039091, -0.040021, -0.009064, 0.025399, -0.029904, -0.018949, -0.025943, -0.003098, -0.003126, -0.035662, -0.006969, -0.112697, -0.109206, -0.193978, -0.182855, -0.191821, -0.241806, -0.210905, -0.251041, -0.167575, -0.107417, -0.016774, 0.007449, 0.019225, 0.008208, -0.028045, 0.005042, -0.046388, -0.021751, -0.036751, -0.018573, -0.030015, 0.032844, 0.005920, -0.025706, 0.002770, -0.019400, -0.013289, -0.048289, -0.146672, -0.176984, -0.222962, -0.207707, -0.271161, -0.249462, -0.216049, -0.191062, -0.160000, -0.082205, -0.040427, -0.050953, -0.014184, 0.008074, 0.017371, -0.011056, -0.080534, -0.060113, -0.036892, 0.016455, -0.031979, 0.012847, -0.009803, 0.012897, 0.010978, -0.021583, -0.002768, -0.061742, -0.169132, -0.140794, -0.148992, -0.161134, -0.190099, -0.159031, -0.168519, -0.144438, -0.096564, -0.086025, -0.068813, -0.091705, -0.001712, -0.031018, -0.000855, -0.026695, -0.056566, -0.021946, 0.002528, 0.029230, -0.005890, 0.034735, 0.009359, 0.020904, -0.008298, 0.022407, 0.013762, -0.096212, -0.077228, -0.137132, -0.123485, -0.115933, -0.056596, -0.061201, -0.028362, -0.031096, -0.023795, -0.090831, -0.060034, -0.042789, -0.021853, -0.049864, -0.030850, -0.084825, -0.095279, -0.053355, -0.032471, 0.035300, -0.015102, -0.002733, 0.014834, -0.031564, 0.027172, -0.015854, -0.012606, -0.047448, -0.052044, -0.042228, -0.038571, 0.018690, 0.030863, 0.095624, 0.104469, 0.104594, 0.036099, 0.021792, 0.041525, 0.019184, -0.047545, -0.035316, -0.075113, -0.042575, -0.056238, 0.006433, 0.015963, 0.027732, -0.012485, -0.026848, 0.005622, -0.017924, -0.017420, 0.031320, 0.002127, 0.010672, 0.065423, 0.053321, 0.026303, 0.079384, 0.110063, 0.091790, 0.152390, 0.125288, 0.063675, 0.091905, 0.043177, 0.058925, -0.010051, -0.032106, 0.020465, -0.007576, 0.014730, 0.046762, 0.017107, 0.020140, 0.029502, 0.032773, -0.003779, 0.025032, 0.011578, 0.024302, 0.026215, 0.112727, 0.109678, 0.091741, 0.108368, 0.064870, 0.120944, 0.130782, 0.157186, 0.143112, 0.110105, 0.101951, 0.057456, 0.033364, 0.034478, 0.022732, 0.012649, 0.091605, 0.077009, 0.059356, 0.107183, 0.078144, -0.003634, 0.018820, -0.022157, 0.012325, 0.031294, 0.040352, 0.084120, 0.105829, 0.134324, 0.137980, 0.118130, 0.110638, 0.146702, 0.143810, 0.149455, 0.115317, 0.082121, 0.064722, 0.113266, 0.068451, 0.018943, 0.036135, 0.080809, 0.086991, 0.109450, 0.122443, 0.107701, 0.058971, 0.009615, 0.023925, 0.022854, 0.029302, -0.004286, -0.002272, 0.068330, 0.091805, 0.153940, 0.140219, 0.127716, 0.114491, 0.161248, 0.165507, 0.163431, 0.095342, 0.083174, 0.057722, 0.025161, 0.027688, 0.074759, 0.050835, 0.123333, 0.142017, 0.159614, 0.164739, 0.117074, 0.059634, 0.026036, -0.014665, -0.018939, -0.006660, 0.017780, 0.038529, 0.089200, 0.090444, 0.127044, 0.118326, 0.166538, 0.118991, 0.103107, 0.125975, 0.068287, 0.020769, -0.005567, -0.012455, 0.049951, 0.008269, 0.107226, 0.137475, 0.132166, 0.148163, 0.176487, 0.138329, 0.111593, 0.054497, -0.019142, 0.022035, 0.018011, -0.025389, 0.016080, -0.008422, 0.018113, 0.069959, 0.089359, 0.099824, 0.090882, 0.135682, 0.120009, 0.046365, -0.004748, -0.012956, -0.063249, -0.061162, -0.013601, 0.063942, 0.058466, 0.112047, 0.104673, 0.098512, 0.112297, 0.090650, 0.044627, 0.040628, 0.016317, 0.022235, 0.013988, 0.003746, 0.018710, -0.017556, 0.039048, 0.048351, 0.028128, 0.053431, 0.033197, 0.025318, 0.034313, 0.014162, -0.031788, -0.049191, -0.106616, -0.091847, -0.011961, -0.027551, 0.060321, 0.102256, 0.111190, 0.097530, 0.042024, 0.053038, 0.009556, -0.004660, 0.027387, -0.012138, -0.025578, -0.028669, 0.022248, 0.000837, 0.034825, 0.004927, -0.043105, -0.015405, -0.008823, -0.033080, -0.054842, -0.102903, -0.117907, -0.093237, -0.141995, -0.099265, -0.082965, -0.034745, -0.007751, -0.014115, 0.007904, 0.059876, 0.028134, 0.031986, -0.012244, 0.030534, -0.007673, -0.012038, 0.007245, -0.012797, -0.014471, -0.007372, -0.007415, -0.033056, -0.014518, -0.079071, -0.042222, -0.047491, -0.083597, -0.097464, -0.119122, -0.068453, -0.048756, -0.041012, -0.056867, -0.033312, 0.002343, -0.019123, -0.032319, -0.040074, 0.013737, 0.013968, 0.034758, -0.016333, 0.015585, -0.011816, -0.008876, 0.020839, -0.032746, 0.025793, 0.014456, -0.026638, 0.007298, -0.029277, -0.026631, -0.043091, -0.068764, -0.036928, -0.014596, -0.034498, -0.044751, -0.022595, -0.016064, -0.030033, -0.045461, -0.034527, -0.016319, 0.005342, 0.027027, -0.001707, 0.012233, 0.020762, -0.015312, -0.011851, 0.023689, 0.025571, 0.008463, -0.027609, 0.020005, -0.030194, 0.016075, 0.000850, 0.007030, -0.039714, -0.018835, 0.007927, 0.020259, -0.017305, 0.025469, -0.013692, -0.027143, -0.020374, -0.001658, -0.009407, 0.014976, -0.020989, -0.010530, -0.035454, 0.029142, -0.006728, -0.028154, -0.001723, -0.000065, 0.009919, -0.003920, 0.022467, -0.012324, -0.010721, -0.008570, 0.006276, 0.028495, -0.001818, 0.027198, 0.027762, -0.019011, -0.003565, -0.017479, 0.014295, -0.013120, 0.010334, 0.001813, -0.023566, -0.024159, -0.034943, -0.020067, 0.009972, 0.002176, 0.026861, -0.031404, -0.001044
--  Sum of weights (converted): 00000000B2284934
    );

    constant weights_n3 : weight_array := (
     x"8106558A", x"0001B66D", x"006A9830", x"81067304", x"0102629C", x"805ADEBB", x"01033A98", x"80311BC2", x"00A5FAEA", x"0109F848", x"806A847B", x"80471EC7", x"009968E4", x"80FADE07", x"00ACE0B9", x"80B7C7D8", x"010FBACA", x"80BFBDBE", x"80786580", x"00DA5003", x"807F61B9", x"00FAC72A", x"00C94B7C", x"010B69E6", x"811B9590", x"00034772", x"80603B10", x"0045B10B", x"80DCE80A", x"0077F857", x"800DDC36", x"808A4B93", x"810732FC", x"0099084B", x"806A0854", x"00D76C10", x"0033512C", x"00581284", x"802D0486", x"8029B9B4", x"80654758", x"80FF5392", x"00B5F194", x"80BA1B09", x"00A8AB43", x"806413CF", x"00B69D8A", x"00FA5B3C", x"80B3534A", x"00F16AAF", x"000718DA", x"80DF8211", x"00776E5C", x"00A5AA5A", x"0101E7B8", x"81168134", x"01082E56", x"00DDCCEE", x"011FD208", x"009F69EA", x"808E609B", x"00DDE50E", x"010AEDB2", x"8071BB65", x"80340CD5", x"00DD01BA", x"00E0F9FA", x"00B8146D", x"00D2E151", x"80AB20DB", x"804A4B16", x"8090160E", x"007FCB80", x"00330EDF", x"80F7F17F", x"80390161", x"80FC8A53", x"811C858A", x"0105346C", x"80952A31", x"00820CF8", x"80412EBA", x"803B3ED9", x"80003060", x"00E42F3E", x"80287922", x"00F21690", x"00AB0B30", x"00C83ED6", x"80FE859A", x"807F917C", x"80E08EFB", x"802A05C9", x"80227282", x"006C60C1", x"0182D12A", x"0148407A", x"00061DEC", x"0032DE7D", x"01A253C2", x"00A86D1C", x"00B6CC2C", x"8062E79A", x"80253FF7", x"003E3B6B", x"80EF847D", x"0098F6CC", x"007D6C25", x"80B3B114", x"80792445", x"8044FFCC", x"002D8822", x"806B5230", x"0117EDCE", x"8119A40A", x"80A2E2A5", x"80A09A2E", x"00947173", x"00AE1DF9", x"00916ADB", x"02645320", x"00E87030", x"02DA07D4", x"02353CC4", x"028E271C", x"0172DDA8", x"00FC5067", x"00220F9E", x"00D1AD19", x"80B446F1", x"002EFD6B", x"8166811C", x"815D3680", x"80F4D6B4", x"0022EE9D", x"80EB7FC4", x"00701995", x"00472E10", x"00B04CF6", x"00B8BFD7", x"0076BAEC", x"80583960", x"80512549", x"0085D847", x"00FF5E57", x"00ED8907", x"024CC454", x"01D44766", x"03F05FF0", x"03C25C9C", x"0383AE5C", x"03AA4120", x"02E5F954", x"036DA374", x"01C1B08C", x"01A61D32", x"01154224", x"80EE1256", x"80BEEFF0", x"8130FCA0", x"810FEEA2", x"810F271A", x"82802C8C", x"80B8443B", x"80A30A69", x"80CB5CEB", x"808A30FA", x"004A4B4C", x"003CEAD4", x"80095DAF", x"808E8B53", x"00D8DB63", x"01178AF0", x"00AE6AD8", x"0292AA9C", x"031E3B58", x"03BC36D8", x"041CB2C0", x"03C1BC78", x"054AE3B8", x"02BAF558", x"04ADE400", x"02A659D8", x"0328A500", x"025B0C94", x"00F1584D", x"015021EC", x"00E7FBDD", x"80AF3D27", x"8175DDB6", x"813F3624", x"81EBE778", x"80B45613", x"00488A60", x"8078BD4D", x"80A387FE", x"006BB175", x"80675EC9", x"80C0CA65", x"802CE865", x"00D6EE81", x"0368FDD0", x"0317FB3C", x"036985F0", x"03141A8C", x"01F1461E", x"02EEB6C0", x"0197A194", x"017DE580", x"02DBDCDC", x"023A630C", x"03C57434", x"02270000", x"02C62B54", x"01CDD4B2", x"00A3EFD8", x"022C6434", x"004F00A5", x"81E151F4", x"80ECCFCD", x"80CC184B", x"800C804A", x"807D8DAF", x"80A16CB3", x"809D6E9D", x"006C8165", x"004703EC", x"804AA0C6", x"026EE390", x"02A17664", x"018F9544", x"01F5CCA8", x"800BAF85", x"801178F0", x"802CA886", x"82AB54FC", x"8206D420", x"809F71D4", x"016CCD06", x"01FCE03A", x"0269BDDC", x"022A2F9C", x"01B1A442", x"026ECE4C", x"027AE6BC", x"01328E92", x"808A58BA", x"81B4231A", x"8158C0AA", x"800EACEF", x"00B71D67", x"80924B29", x"8097EBC5", x"007D9575", x"80DB674F", x"010A2D74", x"01717B60", x"012194B4", x"000CCFBD", x"80AA9E33", x"83418AD0", x"84E9CC40", x"840D77F8", x"86BCEEF0", x"85A58508", x"82C9CB78", x"00E6A621", x"03A1ECB0", x"03355DE8", x"02A415F4", x"01EC3972", x"0349D6E4", x"035B9190", x"016B4E96", x"8072E9C5", x"80791CBD", x"81D76B32", x"002FF9C3", x"80B508FB", x"00E39F91", x"81032DCE", x"0068105C", x"80FABB16", x"00E6D5E5", x"0083912C", x"00D918E6", x"820CA1D0", x"824343A4", x"85BAE850", x"874A6498", x"876A5708", x"87AC55B8", x"85E58510", x"81C463DE", x"0277FF78", x"04EE40B8", x"05914BE0", x"044D7768", x"02B81A44", x"01906CD2", x"009401FD", x"012C688A", x"8172E45E", x"8124B266", x"816FA418", x"80ED5EED", x"00321DEE", x"80488059", x"00212DFB", x"80073239", x"0003BA74", x"8020EC0B", x"801708DA", x"806B9C05", x"8188E874", x"83733BD4", x"870F2A70", x"87E94F30", x"871B0C70", x"853BAD60", x"810F66CA", x"03233894", x"04E62AE8", x"04A26200", x"04976898", x"046214E8", x"02E49F5C", x"0095E6C9", x"001FDA2A", x"8252E134", x"81C68B9E", x"8015864E", x"80DCFFA2", x"00A5C189", x"80F1EABB", x"01029C1C", x"008B79D2", x"00BA1AB3", x"0041F514", x"0003D896", x"80D3D0CA", x"81CDC522", x"837686A8", x"83661EDC", x"85B52710", x"8501BE68", x"84CABB20", x"81126690", x"0197A1E6", x"03861E88", x"05BFCD80", x"041BC350", x"0443F8D0", x"02063360", x"021A3660", x"81397A38", x"8167CCF4", x"81820B4E", x"82776C9C", x"802DF12E", x"00995241", x"80B8434C", x"001727DC", x"00587A44", x"00F24B1F", x"00E286C3", x"80FD2B3A", x"80FA373E", x"814F4844", x"81A2D5EC", x"8295CED4", x"841296E8", x"833E9BC0", x"843BCCD0", x"82E037C0", x"000D62DA", x"035D1DC4", x"0606F3D8", x"0456FA08", x"02F66BD4", x"02F7BF08", x"01AAA3FC", x"00AA6A27", x"80450232", x"80EBFE9B", x"80E5153E", x"816E5428", x"819399E8", x"810FA312", x"0111F55A", x"8109D4A4", x"00448594", x"801C4441", x"011151CA", x"00A92687", x"804A533D", x"81208022", x"80C590A3", x"82E4FFF8", x"83365B28", x"83003B0C", x"82550058", x"81E692BC", x"002BA5FD", x"025818E8", x"01B81DB2", x"01E994DE", x"007F6740", x"01B7A15C", x"0192B7E4", x"00FFEB81", x"0145CB00", x"0074DEED", x"0058B9C7", x"00231522", x"81AAD572", x"8109BD1C", x"80F0E5CE", x"00BFFB97", x"00ABF1B2", x"00ECF455", x"80C81FDC", x"80921805", x"013A37C0", x"80CE72FC", x"814DEB86", x"8136CA26", x"83BEA790", x"83E73544", x"832FFC4C", x"81C27D38", x"80CDCC40", x"807C7B39", x"008F1802", x"00250B31", x"81BA0E88", x"000D25A1", x"00A9AC1E", x"01CD4DA6", x"029FB5DC", x"02692E18", x"01790F74", x"80F9ACCD", x"80BF99B9", x"0019DB9A", x"803C39C0", x"805F2D4E", x"8097B450", x"011561B2", x"80E62E47", x"80C0DA63", x"0141EF36", x"8015B621", x"00A399D5", x"81E524DA", x"8299140C", x"84692E10", x"83C579E0", x"8414AAB0", x"83E258BC", x"8354F69C", x"84189178", x"84AF8B88", x"838A09F8", x"80731B4E", x"015DC8F8", x"03E82598", x"035EFD64", x"02BCAF30", x"01770788", x"0156A022", x"812C08A8", x"801649FC", x"003A629F", x"002C2759", x"00CD05E9", x"00463815", x"804EA4A1", x"809711CF", x"802F41EB", x"01E089F8", x"012C37C6", x"81A9E53E", x"81C71078", x"843457A0", x"84BE8F98", x"8705D160", x"85B0A130", x"857B7730", x"85CC7F40", x"857396D8", x"837B63EC", x"0002C349", x"0192FB24", x"032CB3E4", x"0380CFD8", x"036745C8", x"02219AD4", x"01E15C1A", x"00D1DED1", x"80187973", x"0054DF19", x"802EF616", x"008B9A88", x"80649678", x"00FED8F6", x"00472A9E", x"016BF8B4", x"0145E890", x"02D69EF4", x"0037DDCC", x"80618C5E", x"83BA8408", x"86174098", x"868C0438", x"87733DF8", x"866D5D10", x"86A295B0", x"866596A0", x"821E5B48", x"01C51564", x"023BB880", x"031E404C", x"04638520", x"0264BDF4", x"02F6A514", x"0110E944", x"8002E268", x"815A91C0", x"803D4CD0", x"806F7DDF", x"80842970", x"808FD7D8", x"00433155", x"0123A7BE", x"01ED20E0", x"03076ED4", x"041037B8", x"02C5EDDC", x"00578684", x"82191278", x"82DDF2C0", x"83FF49A4", x"85D50950", x"860ABF40", x"847EB240", x"825D4E18", x"81FCAF7E", x"0153E79C", x"03579EE4", x"0318AAD4", x"031274CC", x"03F9F148", x"03303B3C", x"801F036E", x"8080718B", x"818A2202", x"0045D8C3", x"80CF5A2A", x"80954DA7", x"80879C2A", x"002D077B", x"01242446", x"0193F700", x"03A9A16C", x"04DF3788", x"03333070", x"0250F4D0", x"013BCFFC", x"806DCCE6", x"814C648A", x"821565A4", x"8378B820", x"812A644A", x"8025162E", x"00A30BE1", x"037D289C", x"0383FDBC", x"0467CC90", x"022D5A34", x"03A7D84C", x"025F5FA4", x"8105C590", x"81B89CA2", x"80D79ECD", x"80D57719", x"0049ED8D", x"008236E1", x"8025498B", x"00CF059E", x"006294D7", x"013ADA48", x"020291F4", x"043D10C0", x"030C7E24", x"03890B18", x"02F7801C", x"00BC26FC", x"00710788", x"80BF77B0", x"8039F15E", x"006D7696", x"80279B05", x"010C8C10", x"023E4A5C", x"01E8A148", x"030D7AA4", x"017C821E", x"00612190", x"0043DEFC", x"800D9606", x"810ADA56", x"81874710", x"00130E36", x"00938E28", x"00E48C33", x"001BC047", x"00CB2FE5", x"80C8E997", x"0216020C", x"016D49C0", x"0235F830", x"04A27E18", x"039B66F0", x"0414D0A8", x"0248A7C4", x"03249098", x"02AF3E60", x"01743476", x"0245F384", x"00BC7FB5", x"0181AF70", x"01DD27B4", x"01FB2A20", x"008A2956", x"0184E874", x"8069E4BE", x"8147C454", x"8067EDA5", x"815245EE", x"813C3988", x"005690EA", x"00636EE3", x"007081A9", x"80265E0D", x"80D5F7C5", x"80D42FC3", x"019F69A0", x"006C4870", x"02986FE8", x"04108660", x"047F2D60", x"02C2128C", x"033437F8", x"0267A01C", x"0395B770", x"0139DD10", x"011A412C", x"0094AC19", x"01997EAA", x"00B2913E", x"00DB961B", x"0124C674", x"80A9AB4D", x"812FEDA2", x"8141DBDE", x"8005AADE", x"003D75AD", x"002CC262", x"80E5767C", x"001A42FA", x"809B4017", x"80398887", x"802D4AF0", x"00136823", x"80CA8BCA", x"01A0AC3A", x"00AF9E55", x"0238E320", x"03402C88", x"034C9E9C", x"03E15FF8", x"03DF9898", x"03E5F138", x"02DA3B08", x"03078ABC", x"00D73BBB", x"80182CD1", x"00A753FF", x"00109CEA", x"809BF820", x"817A63B2", x"800C0F30", x"007AF95C", x"80489119", x"0030201C", x"00797C89", x"8122F058", x"80302B03", x"806C88A5", x"809589E5", x"00B2D275", x"01228A12", x"002FC76B", x"00CAC888", x"80A89191", x"008CE141", x"005C6B83", x"00143859", x"012FDC00", x"0179C9D2", x"011EE18C", x"01B90A52", x"0183D73C", x"01865C86", x"001794DE", x"80351DF2", x"80762171", x"803236E7", x"80E8B326", x"8048A69A", x"810FB9DC", x"80D78C6E", x"80FED1BC", x"00D77DD2", x"80A838FC", x"80179E01", x"001F4749", x"0102676A", x"0084C7D5", x"80D0598E", x"011E1E00", x"8115C288", x"00266FEE", x"01090414", x"00F987F7", x"805598AE", x"80E21236", x"004E6AD2", x"00A2F622", x"80E090F5", x"80766F21", x"810955D4", x"00185D25", x"80109FE8", x"00505775", x"808A9512", x"812C1480", x"8083908C", x"80E96A79", x"80479E03", x"0069E77B", x"80F379CF", x"800DAB97", x"811E3F00", x"80CF54A1", x"80CCD731", x"80639DC5", x"80943D4E", x"002D08A9", x"00B2D842", x"00DC6322", x"005BA22A", x"80029A66", x"80356C27", x"00C45889", x"80AB73B6", x"00CF42BC", x"81203474", x"80E435C9", x"003F6CE9", x"80863639", x"00266350", x"00F032F7", x"007C70EE", x"011A17EE", x"807DAF4A", x"808C5FCD", x"80259D77", x"803AF780", x"8080B17E", x"80122A26", x"0108509C", x"80A06013"
--  -0.032023, 0.000209, 0.013012, -0.032037, 0.031541, -0.011093, 0.031644, -0.005995, 0.020261, 0.032467, -0.013003, -0.008682, 0.018727, -0.030623, 0.021103, -0.022434, 0.033170, -0.023406, -0.014697, 0.026649, -0.015550, 0.030613, 0.024572, 0.032643, -0.034617, 0.000400, -0.011747, 0.008507, -0.026966, 0.014645, -0.001692, -0.016882, -0.032129, 0.018681, -0.012943, 0.026297, 0.006264, 0.010751, -0.005495, -0.005093, -0.012363, -0.031168, 0.022210, -0.022718, 0.020589, -0.012216, 0.022292, 0.030561, -0.021890, 0.029470, 0.000866, -0.027284, 0.014579, 0.020223, 0.031483, -0.033997, 0.032249, 0.027075, 0.035134, 0.019460, -0.017380, 0.027087, 0.032584, -0.013883, -0.006354, 0.026978, 0.027463, 0.022471, 0.025742, -0.020890, -0.009069, -0.017589, 0.015600, 0.006233, -0.030267, -0.006959, -0.030828, -0.034732, 0.031885, -0.018209, 0.015875, -0.007957, -0.007232, -0.000023, 0.027855, -0.004941, 0.029552, 0.020879, 0.024444, -0.031070, -0.015572, -0.027412, -0.005130, -0.004205, 0.013230, 0.047219, 0.040070, 0.000747, 0.006210, 0.051065, 0.020560, 0.022314, -0.012073, -0.004547, 0.007597, -0.029238, 0.018672, 0.015310, -0.021935, -0.014788, -0.008423, 0.005558, -0.013101, 0.034171, -0.034380, -0.019883, -0.019605, 0.018121, 0.021255, 0.017751, 0.074747, 0.028374, 0.089115, 0.068999, 0.079853, 0.045272, 0.030800, 0.004158, 0.025595, -0.022006, 0.005736, -0.043763, -0.042629, -0.029888, 0.004264, -0.028747, 0.013684, 0.008689, 0.021521, 0.022552, 0.014493, -0.010770, -0.009905, 0.016338, 0.031173, 0.028996, 0.071871, 0.057163, 0.123093, 0.117476, 0.109824, 0.114533, 0.090573, 0.107134, 0.054894, 0.051528, 0.033845, -0.029061, -0.023308, -0.037230, -0.033195, -0.033100, -0.078146, -0.022493, -0.019902, -0.024825, -0.016869, 0.009069, 0.007436, -0.001143, -0.017400, 0.026472, 0.034124, 0.021291, 0.080404, 0.097440, 0.116725, 0.128503, 0.117399, 0.165392, 0.085322, 0.146227, 0.082807, 0.098711, 0.073614, 0.029461, 0.041032, 0.028318, -0.021391, -0.045638, -0.038966, -0.060047, -0.022014, 0.008855, -0.014739, -0.019962, 0.013146, -0.012618, -0.023534, -0.005482, 0.026237, 0.106566, 0.096677, 0.106631, 0.096204, 0.060702, 0.091640, 0.049760, 0.046618, 0.089339, 0.069627, 0.117853, 0.067261, 0.086691, 0.056376, 0.020012, 0.067919, 0.009644, -0.058755, -0.028908, -0.024914, -0.001526, -0.015326, -0.019705, -0.019218, 0.013245, 0.008669, -0.009110, 0.076036, 0.082210, 0.048777, 0.061255, -0.001426, -0.002133, -0.005451, -0.083415, -0.063334, -0.019463, 0.044531, 0.062119, 0.075408, 0.067650, 0.052935, 0.076026, 0.077503, 0.037421, -0.016888, -0.053239, -0.042084, -0.001791, 0.022353, -0.017858, -0.018545, 0.015330, -0.026783, 0.032492, 0.045103, 0.035349, 0.001564, -0.020827, -0.101751, -0.153540, -0.126644, -0.210563, -0.176455, -0.087133, 0.028155, 0.113516, 0.100265, 0.082530, 0.060086, 0.102764, 0.104928, 0.044349, -0.014027, -0.014784, -0.057546, 0.005856, -0.022099, 0.027786, -0.031638, 0.012703, -0.030607, 0.028178, 0.016060, 0.026501, -0.064042, -0.070711, -0.179066, -0.227831, -0.231731, -0.239787, -0.184268, -0.055223, 0.077148, 0.154084, 0.173986, 0.134456, 0.084973, 0.048880, 0.018067, 0.036671, -0.045275, -0.035730, -0.044878, -0.028976, 0.006118, -0.008850, 0.004050, -0.000878, 0.000455, -0.004019, -0.002812, -0.013136, -0.047962, -0.107817, -0.220601, -0.247230, -0.222052, -0.163535, -0.033130, 0.098049, 0.153097, 0.144822, 0.143482, 0.136973, 0.090408, 0.018299, 0.003888, -0.072617, -0.055486, -0.002628, -0.026977, 0.020234, -0.029531, 0.031569, 0.017026, 0.022718, 0.008051, 0.000469, -0.025856, -0.056368, -0.108219, -0.106216, -0.178363, -0.156463, -0.149747, -0.033496, 0.049760, 0.110122, 0.179663, 0.128389, 0.133297, 0.063257, 0.065700, -0.038266, -0.043921, -0.047125, -0.077078, -0.005608, 0.018716, -0.022493, 0.002827, 0.010800, 0.029577, 0.027652, -0.030904, -0.030544, -0.040928, -0.051127, -0.080787, -0.127269, -0.101393, -0.132300, -0.089870, 0.001634, 0.105117, 0.188349, 0.135617, 0.092581, 0.092742, 0.052080, 0.020803, -0.008424, -0.028808, -0.027964, -0.044718, -0.049268, -0.033159, 0.033442, -0.032450, 0.008364, -0.003451, 0.033364, 0.020648, -0.009073, -0.035217, -0.024117, -0.090454, -0.100385, -0.093778, -0.072876, -0.059396, 0.005328, 0.073254, 0.053725, 0.059763, 0.015552, 0.053666, 0.049160, 0.031240, 0.039770, 0.014266, 0.010831, 0.004283, -0.052104, -0.032439, -0.029406, 0.023435, 0.020989, 0.028925, -0.024429, -0.017834, 0.038357, -0.025201, -0.040762, -0.037938, -0.117023, -0.121974, -0.099608, -0.054991, -0.025122, -0.015195, 0.017468, 0.004522, -0.053962, 0.001605, 0.020712, 0.056311, 0.081996, 0.075339, 0.046028, -0.030478, -0.023389, 0.003156, -0.007352, -0.011618, -0.018519, 0.033860, -0.028098, -0.023542, 0.039299, -0.002650, 0.019971, -0.059222, -0.081186, -0.137839, -0.117856, -0.127523, -0.121380, -0.104121, -0.127999, -0.146429, -0.110600, -0.014051, 0.042698, 0.122088, 0.105345, 0.085533, 0.045780, 0.041824, -0.036625, -0.002721, 0.007127, 0.005390, 0.025027, 0.008572, -0.009600, -0.018441, -0.005769, 0.058660, 0.036648, -0.051989, -0.055550, -0.131389, -0.148262, -0.219460, -0.177811, -0.171321, -0.181213, -0.170360, -0.108812, 0.000337, 0.049192, 0.099207, 0.109474, 0.106357, 0.066602, 0.058760, 0.025619, -0.002988, 0.010360, -0.005733, 0.017041, -0.012279, 0.031109, 0.008687, 0.044430, 0.039784, 0.088699, 0.006820, -0.011908, -0.116518, -0.190338, -0.204592, -0.232818, -0.200850, -0.207347, -0.199901, -0.066206, 0.055308, 0.069790, 0.097443, 0.137148, 0.074798, 0.092608, 0.033314, -0.000352, -0.042306, -0.007483, -0.013610, -0.016133, -0.017559, 0.008202, 0.035602, 0.060196, 0.094657, 0.126980, 0.086661, 0.010684, -0.065561, -0.089593, -0.124913, -0.182255, -0.188812, -0.140466, -0.073890, -0.062095, 0.041492, 0.104446, 0.096761, 0.096003, 0.124261, 0.099638, -0.003786, -0.015679, -0.048112, 0.008526, -0.025312, -0.018226, -0.016554, 0.005497, 0.035662, 0.049312, 0.114457, 0.152248, 0.099999, 0.072382, 0.038551, -0.013403, -0.040575, -0.065112, -0.108486, -0.036425, -0.004527, 0.019903, 0.109028, 0.109862, 0.137671, 0.068036, 0.114239, 0.074142, -0.031955, -0.053786, -0.026321, -0.026058, 0.009024, 0.015895, -0.004552, 0.025271, 0.012034, 0.038434, 0.062814, 0.132454, 0.095275, 0.110479, 0.092712, 0.022968, 0.013798, -0.023373, -0.007073, 0.013362, -0.004835, 0.032782, 0.070104, 0.059647, 0.095395, 0.046449, 0.011857, 0.008285, -0.001658, -0.032575, -0.047763, 0.002326, 0.018012, 0.027899, 0.003388, 0.024803, -0.024525, 0.065187, 0.044591, 0.069088, 0.144836, 0.112720, 0.127541, 0.071369, 0.098213, 0.083892, 0.045435, 0.071039, 0.023010, 0.047081, 0.058246, 0.061910, 0.016865, 0.047474, -0.012926, -0.040011, -0.012687, -0.041293, -0.038602, 0.010567, 0.012138, 0.013734, -0.004684, -0.026119, -0.025902, 0.050710, 0.013218, 0.081108, 0.127017, 0.140525, 0.086190, 0.100124, 0.075150, 0.112026, 0.038313, 0.034455, 0.018148, 0.049987, 0.021798, 0.026805, 0.035739, -0.020712, -0.037101, -0.039289, -0.000692, 0.007502, 0.005464, -0.028011, 0.003206, -0.018951, -0.007023, -0.005529, 0.002369, -0.024725, 0.050863, 0.021438, 0.069444, 0.101584, 0.103103, 0.121262, 0.121044, 0.121819, 0.089139, 0.094671, 0.026274, -0.002951, 0.020426, 0.002028, -0.019039, -0.046190, -0.001472, 0.015011, -0.008858, 0.005875, 0.014830, -0.035515, -0.005880, -0.013249, -0.018254, 0.021829, 0.035466, 0.005832, 0.024754, -0.020577, 0.017197, 0.011282, 0.002468, 0.037092, 0.046117, 0.035020, 0.053838, 0.047344, 0.047652, 0.002879, -0.006484, -0.014420, -0.006130, -0.028406, -0.008869, -0.033170, -0.026312, -0.031106, 0.026305, -0.020535, -0.002883, 0.003818, 0.031543, 0.016209, -0.025433, 0.034926, -0.033906, 0.004692, 0.032351, 0.030460, -0.010449, -0.027597, 0.009572, 0.019893, -0.027413, -0.014457, -0.032390, 0.002974, -0.002029, 0.009807, -0.016917, -0.036631, -0.016060, -0.028493, -0.008742, 0.012928, -0.029721, -0.001669, -0.034942, -0.025309, -0.025005, -0.012160, -0.018096, 0.005497, 0.021832, 0.026903, 0.011186, -0.000318, -0.006521, 0.023968, -0.020929, 0.025300, -0.035181, -0.027858, 0.007742, -0.016383, 0.004686, 0.029321, 0.015191, 0.034435, -0.015342, -0.017136, -0.004592, -0.007198, -0.015710, -0.002217, 0.032265, -0.019577
--  Sum of weights (converted): 00000000856AE45C
    );

    constant weights_n4 : weight_array := (
     x"00A44D9A", x"0087E9AE", x"00A96EF0", x"004EEE27", x"806C148E", x"0078BF89", x"8089CCC5", x"80B395DC", x"01117E8C", x"00F28243", x"80D3713E", x"00EDA465", x"003BC2EF", x"0048327E", x"0119187C", x"800F6665", x"805D0D45", x"00B7AB53", x"804B9345", x"80463C35", x"8075FB20", x"011FF98C", x"008B9A83", x"802F6DD7", x"8005D640", x"001479F6", x"80AD6F71", x"00531177", x"80E312B1", x"800DA424", x"8036E589", x"80777635", x"010E91F8", x"0051D221", x"0089BA6F", x"80C7E4FD", x"00243D76", x"0043A248", x"0083EAF0", x"807226EF", x"805C0828", x"81056956", x"00A36181", x"00B2B135", x"00764706", x"008932D8", x"00A87407", x"010F0406", x"005BCB14", x"00666C0D", x"0059A87C", x"80A640A8", x"004967D0", x"0058263E", x"80E8DF81", x"80569697", x"80B483D5", x"80BAF0F1", x"00CB5140", x"00E61395", x"80297CDC", x"00593B0B", x"80499D20", x"0027F128", x"8056947D", x"80D344B2", x"80E3B37D", x"00904907", x"80828124", x"814BA3FC", x"807D32AF", x"81B53B72", x"807CA5EF", x"007D18BC", x"80280074", x"001B3CD0", x"812CF62E", x"804C0CFF", x"009EC996", x"80DCEFC8", x"808BBB52", x"00C4AC9E", x"00540530", x"0088C4F5", x"8110D3EE", x"00BA34F7", x"803FD338", x"003D04E1", x"00EBAF3B", x"81103A4C", x"0046BFB8", x"812ED4E6", x"00887343", x"80391DCC", x"80BF4875", x"81A544CC", x"8105C20E", x"8231DEE0", x"81616C5C", x"80972C67", x"8239B51C", x"817909F0", x"8093EF54", x"80518534", x"80411930", x"00D4352C", x"8062CC80", x"0045B2A6", x"009478EC", x"803A5D40", x"00BEE67E", x"00BF140E", x"0082482E", x"80476167", x"00FE15DC", x"80A97C41", x"005D5EB7", x"003DD509", x"00C1711B", x"8115657E", x"8036E206", x"817CB226", x"80D4668E", x"816561EA", x"83110B48", x"828DAE44", x"82672608", x"8225A480", x"8119D6E4", x"81146E0A", x"80E9C419", x"000E6CC1", x"80F3934B", x"011696D8", x"004964A1", x"010A0910", x"0086EE55", x"8008F196", x"00CD5BEA", x"80AADA6B", x"0052816E", x"00804195", x"806837A7", x"0069D447", x"8117C5A6", x"80778AC2", x"00C7BC5C", x"00CB73D8", x"8111AC66", x"00127384", x"80EE8772", x"807B46BE", x"832CFBA8", x"82ED21E0", x"837A4154", x"834B9EA8", x"81B37706", x"81981096", x"0145149A", x"0089A82A", x"01C23EB6", x"00FC4B4A", x"01D4D2B8", x"00E77C48", x"01AC8134", x"010EAB60", x"00E088AE", x"8066A56D", x"00B617BA", x"80F47213", x"0084DFAE", x"80286AEA", x"80DF94BC", x"80AB633A", x"80AD4ACF", x"00C52382", x"802B5392", x"80C5ECC0", x"0003F9C8", x"8280ABF0", x"82C98AC0", x"84E59BF0", x"859FD348", x"8633BBF8", x"8443AD20", x"828A6818", x"8143D3FC", x"01538DC4", x"0145CF98", x"01A75AFE", x"032F31A0", x"026176B0", x"002F377E", x"0043B211", x"80445F7F", x"80763347", x"808BA2EB", x"807CBB4E", x"8079E577", x"0013CF21", x"01216A88", x"807590B8", x"80548BD3", x"809A8361", x"80447C25", x"809B4D98", x"827F822C", x"82C071E0", x"85EFD770", x"85DC8640", x"8923AFE0", x"8A1B88D0", x"883EB040", x"84063820", x"8170D1B2", x"81ABD7E2", x"0002E71E", x"0289E650", x"020C3284", x"00EE7F2D", x"001406AA", x"8013FFFE", x"804482E2", x"80CA01A0", x"80B767C3", x"004BA6C1", x"00B9B79D", x"00E8D618", x"80374AD0", x"006E2AFF", x"812A4210", x"00252E0E", x"002D6A3B", x"80842DE5", x"8299D6C4", x"822E5984", x"856861F0", x"86349AC0", x"89166B70", x"8A65B880", x"87204848", x"83DE0224", x"81152F30", x"80E8ECCF", x"0070EFF3", x"0094529C", x"01CBCF0E", x"00836C74", x"009F4F2C", x"007A0FDC", x"811CF024", x"80C72EE3", x"00AF76B5", x"010EBB18", x"811289B4", x"803F8C8F", x"80BD56F7", x"00BC5616", x"00333ECD", x"000812DD", x"804DEA9C", x"8124C080", x"80363208", x"81B3ABE8", x"8187014A", x"841E90A8", x"87F838D8", x"872F63F0", x"829F40EC", x"80345042", x"807F387C", x"80651572", x"80284838", x"80E0EDEA", x"004B9472", x"81B259AA", x"80F55B41", x"8188F5EE", x"81309C2E", x"80283F92", x"0108685C", x"010E427A", x"004BF0FC", x"0098E883", x"81005690", x"0011E725", x"803A8AB5", x"81BDDDE4", x"811ACC20", x"00E305BA", x"01316548", x"00F7AE80", x"00411ABE", x"81D92F1A", x"85C1D268", x"840D9C40", x"81209B72", x"0374B308", x"00858088", x"00835196", x"80D0EA05", x"80EA13CD", x"809120DF", x"8174BF30", x"811F8FB6", x"0076AC20", x"80FE91BC", x"008063F3", x"804BF365", x"8068A30C", x"00A1CF69", x"8007BC4E", x"816E057C", x"0081D135", x"80FEC876", x"012A3C82", x"00E9374C", x"03A85D04", x"047E9AE0", x"047335F8", x"027393CC", x"82FE51EC", x"858CCC98", x"816B7D48", x"03787A18", x"03F0A90C", x"02E60088", x"800CAE95", x"81E3F47E", x"82015690", x"809CF131", x"8195060E", x"001CB0CF", x"815748CA", x"8001D95E", x"80CAA473", x"0067B04A", x"00E7BDCB", x"005960D4", x"8093C887", x"81652AFE", x"80B46631", x"001D9F6F", x"0327B828", x"02F12E2C", x"057E1AA8", x"07B911F8", x"065B5980", x"011761CA", x"828AB110", x"841727B8", x"0023AA6B", x"04020918", x"04B17470", x"030211E8", x"002FDAD6", x"80967AF9", x"815BB460", x"80422CF2", x"80A81A4A", x"808854F2", x"00280039", x"80EE74C8", x"00098E98", x"00862CF5", x"81143770", x"80AB0930", x"009530D3", x"0006DB98", x"00A88717", x"02AD6D9C", x"03D00FA0", x"067BB4D0", x"06E4CE28", x"07D9D668", x"0740DE58", x"016B806C", x"816804CA", x"81EA126C", x"006F816C", x"057E9588", x"04C21630", x"02CA605C", x"00ADA6F8", x"01AAA64C", x"0080EDC8", x"812894C4", x"80020B1D", x"804CF636", x"0100D970", x"009E0018", x"80ADB842", x"0104C5EA", x"80355402", x"8048E8C6", x"0056A7A7", x"01A57DD4", x"0223AF6C", x"03134ED0", x"05C37DA0", x"080DA890", x"07404CD8", x"0759F6A0", x"0560C450", x"02C7BD38", x"8008C84A", x"002239FC", x"0313DFC4", x"07744698", x"07CC3A10", x"04D6E140", x"042A2120", x"0304B78C", x"0015AA78", x"00D4D5FC", x"80DE280D", x"00AA59DD", x"80952577", x"0033ABA3", x"800366C0", x"0087B6D7", x"002D6913", x"80D37EA4", x"008B25DB", x"0149B38A", x"0194619A", x"03C97BE0", x"05918818", x"06ABFD78", x"06AC8380", x"063E1800", x"055DE6B8", x"0384B340", x"02DF6880", x"02DDD008", x"05083430", x"07DFE3C0", x"06F5E608", x"050A8980", x"03077878", x"0293CF3C", x"002B7E74", x"00B545BC", x"00B0C0DD", x"813290E0", x"80C7C8B5", x"80EC0BCA", x"004D7654", x"00388659", x"809717C4", x"00AE5166", x"006EDE15", x"80D61090", x"0180B5C6", x"03231570", x"04FAEB08", x"066F8AC0", x"04D97DF0", x"03243E1C", x"044D9F70", x"02607A94", x"031AB0B4", x"05AB9E80", x"08BCF5F0", x"09626EA0", x"0644C530", x"04C88910", x"019744B2", x"01054BAC", x"802E363A", x"802E2D10", x"814AE6AE", x"802DC5DD", x"00585A7A", x"00D27518", x"803276F8", x"010B4B8C", x"8114788A", x"80533477", x"002B4E75", x"80065CA4", x"00D74DD4", x"00BC8167", x"033BECCC", x"01BE3208", x"014D51D2", x"012D8424", x"00235D59", x"010FBBA4", x"02D3749C", x"06A38F88", x"0713C978", x"05B323E8", x"03613BA4", x"0093852B", x"813FA642", x"81D426BC", x"826F52F8", x"80BED1C3", x"81689B18", x"80EA3A23", x"81418C06", x"0022233B", x"802D72DA", x"80C798B9", x"00BB87D3", x"00F42CC6", x"8123762E", x"801D3FD8", x"810C301E", x"80DE66D2", x"80380EDE", x"81120D0C", x"80B55F37", x"81EB32D6", x"82D6BBC4", x"80B9F86F", x"00F4C259", x"03C1C814", x"02E2CE34", x"01AC53EC", x"80994C90", x"8294B024", x"834394B0", x"81803D20", x"81B79B44", x"80FCD972", x"81B897A4", x"810B8C5C", x"809D6B6B", x"0002FE61", x"80D22618", x"002AE434", x"80BC381E", x"0029C8B9", x"00C6DC1B", x"80AC07FF", x"80B67C81", x"83446CDC", x"837AD8C4", x"84E77CD0", x"8517FE00", x"85C76818", x"8504BF90", x"83A1817C", x"80C0BF59", x"00BB6335", x"0092F021", x"80FEE217", x"80644E12", x"8173D30E", x"8380CB9C", x"829D81D8", x"81756F1C", x"82D6F6A8", x"81ED03B2", x"0033A648", x"802A94F7", x"005ACCB6", x"8079AE88", x"00350BD9", x"00C1CE2A", x"804B63BA", x"809CC429", x"81E3FD50", x"81D9C08A", x"822C2B28", x"854EB638", x"85824660", x"854B90C0", x"86681448", x"85469600", x"83A2E73C", x"82C2BA5C", x"81906E24", x"823CB028", x"808A7E22", x"81909902", x"82097654", x"8254CCE0", x"816343A6", x"82409280", x"82229040", x"8167928C", x"8115C10A", x"80A51316", x"00E51DEF", x"80E257EE", x"80ABFB86", x"80EE8724", x"809737F9", x"8036642D", x"813CFBF8", x"813FA4D6", x"821F0700", x"83F0230C", x"84301D98", x"84F83318", x"83EF80C4", x"84127C88", x"8240E3D8", x"8229102C", x"820AE870", x"80F5B05C", x"81CB45E4", x"815A3FD8", x"802E5D42", x"8070A031", x"002A5673", x"80CEC729", x"80B45B9A", x"008299BD", x"801B9889", x"01022F7A", x"8096F50A", x"805FFE48", x"000CA3FE", x"009C0A40", x"8102C6EA", x"806D2ABA", x"00807558", x"8099F358", x"80DAEFD0", x"82F75BB0", x"84033FC0", x"846FFA80", x"84040030", x"83A81888", x"81FE9256", x"822C4754", x"82D99948", x"0032D124", x"00342102", x"01205338", x"00515E01", x"0167982A", x"8081F7FB", x"00FF98DE", x"80B53B06", x"005D9B1D", x"80772005", x"00B6F7D5", x"80F571E9", x"80390B94", x"804EF845", x"80AEF315", x"80906DF9", x"805B9D02", x"800C62A3", x"00552DF5", x"811A6018", x"804987CC", x"82569F8C", x"828CD3E0", x"81F7EAF4", x"81E0F616", x"818452EE", x"80DFE511", x"80EBBE43", x"81072778", x"00491738", x"014A36FE", x"00B29CEB", x"01A1E03C", x"01ECF26E", x"01006676", x"0007326E", x"801F7A98", x"80910166", x"8021D220", x"0100C326", x"80966AE3", x"002ECEA7", x"80D6AA7C", x"80502242", x"000E6A81", x"80EFF726", x"001B007C", x"8162B6E6", x"811F2A7C", x"80122800", x"0006B239", x"813FB3D0", x"81E0FBD0", x"826BE3F8", x"81FB9F5A", x"81CD6164", x"00337649", x"810B4EDA", x"00C90273", x"00BBB604", x"00077A94", x"011153E4", x"00A50F16", x"80162EF9", x"80D5796D", x"805E5385", x"005EE576", x"00FD69EF", x"8062BB07", x"80799677", x"811DDB6E", x"00B3C32C", x"011D2662", x"00C472BA", x"80BBEF42", x"00928D43", x"80E3705B", x"805621F4", x"8099FDE6", x"82983278", x"81FD252A", x"822C7464", x"834AF338", x"8171B0D6", x"817C3A5E", x"81617CF8", x"8229FCD0", x"8234DAA4", x"81CF4166", x"8062F1A4", x"80B72E3E", x"00B58792", x"00E50756", x"000FFBA7", x"80F01D09", x"00740A06", x"0105D21C", x"80497C29", x"80991E17", x"804470B7", x"0029DEC5", x"80DB676C", x"0095A3E3", x"006151AE", x"80AE4CE6", x"80E1638C", x"81393752", x"00003CDD", x"8081E4C9", x"8104C84C", x"817F0114", x"81450788", x"8047CAE2", x"80F4246F", x"81A97F6C", x"8066703D", x"810A504C", x"80631865", x"80E7180E", x"80171AEE", x"000DFD9C", x"80B17D34", x"00BC0D1D", x"010E3738", x"80F4B7AA", x"0054C6DE", x"80CA1C05", x"803A269B", x"008C2580", x"80052732", x"00580E78", x"806116CA", x"010F1CFA", x"8093B7A9", x"002C5B70", x"000CA5D6", x"00B4C019", x"000647A9", x"0093B5A0", x"001CC110", x"0097C294", x"801E6AC7", x"00420BF4", x"0107410E", x"806E9F2F", x"807D3556", x"00D0FBCF", x"006CC537", x"8114785C", x"00680E89", x"811EF0D0", x"809ED7FC", x"00727EFE"
--  0.020057, 0.016591, 0.020683, 0.009635, -0.013193, 0.014740, -0.016821, -0.021922, 0.033386, 0.029603, -0.025811, 0.029009, 0.007295, 0.008813, 0.034313, -0.001880, -0.011359, 0.022421, -0.009225, -0.008574, -0.014402, 0.035153, 0.017041, -0.005790, -0.000713, 0.002500, -0.021171, 0.010140, -0.027719, -0.001665, -0.006701, -0.014583, 0.033029, 0.009988, 0.016813, -0.024401, 0.004424, 0.008256, 0.016103, -0.013935, -0.011234, -0.031911, 0.019944, 0.021813, 0.014438, 0.016748, 0.020563, 0.033083, 0.011205, 0.012503, 0.010945, -0.020295, 0.008961, 0.010760, -0.028427, -0.010570, -0.022036, -0.022820, 0.024819, 0.028086, -0.005064, 0.010892, -0.008986, 0.004876, -0.010569, -0.025790, -0.027796, 0.017613, -0.015931, -0.040483, -0.015283, -0.053373, -0.015216, 0.015271, -0.004883, 0.003325, -0.036738, -0.009284, 0.019383, -0.026970, -0.017057, 0.024008, 0.010256, 0.016695, -0.033304, 0.022730, -0.007791, 0.007449, 0.028770, -0.033231, 0.008636, -0.036967, 0.016657, -0.006972, -0.023350, -0.051424, -0.031953, -0.068588, -0.043142, -0.018454, -0.069544, -0.046025, -0.018058, -0.009951, -0.007947, 0.025904, -0.012060, 0.008508, 0.018124, -0.007125, 0.023303, 0.023325, 0.015904, -0.008713, 0.031016, -0.020689, 0.011398, 0.007548, 0.023614, -0.033862, -0.006700, -0.046472, -0.025928, -0.043626, -0.095831, -0.079795, -0.075091, -0.067095, -0.034404, -0.033744, -0.028536, 0.001761, -0.029733, 0.034007, 0.008959, 0.032475, 0.016471, -0.001092, 0.025068, -0.020856, 0.010071, 0.015656, -0.012722, 0.012919, -0.034152, -0.014593, 0.024382, 0.024836, -0.033407, 0.002252, -0.029117, -0.015048, -0.099241, -0.091447, -0.108674, -0.102981, -0.053157, -0.049813, 0.039683, 0.016804, 0.054962, 0.030798, 0.057229, 0.028258, 0.052308, 0.033041, 0.027409, -0.012530, 0.022228, -0.029840, 0.016220, -0.004934, -0.027293, -0.020921, -0.021154, 0.024065, -0.005289, -0.024161, 0.000485, -0.078207, -0.087102, -0.153028, -0.175760, -0.193815, -0.133261, -0.079395, -0.039530, 0.041449, 0.039772, 0.051679, 0.099511, 0.074397, 0.005764, 0.008264, -0.008346, -0.014429, -0.017045, -0.015226, -0.014880, 0.002418, 0.035329, -0.014351, -0.010321, -0.018861, -0.008360, -0.018958, -0.078065, -0.085992, -0.185528, -0.183169, -0.285606, -0.315861, -0.257652, -0.125759, -0.045022, -0.052227, 0.000354, 0.079333, 0.063989, 0.029113, 0.002445, -0.002441, -0.008363, -0.024659, -0.022388, 0.009235, 0.022671, 0.028422, -0.006750, 0.013448, -0.036408, 0.004539, 0.005544, -0.016135, -0.081279, -0.068158, -0.168992, -0.193921, -0.283987, -0.324917, -0.222691, -0.120851, -0.033836, -0.028433, 0.013786, 0.018106, 0.056129, 0.016043, 0.019447, 0.014900, -0.034782, -0.024314, 0.021419, 0.033048, -0.033513, -0.007757, -0.023113, 0.022990, 0.006256, 0.000986, -0.009511, -0.035736, -0.006616, -0.053183, -0.047730, -0.128731, -0.249051, -0.224535, -0.081940, -0.006386, -0.015530, -0.012339, -0.004917, -0.027457, 0.009226, -0.053021, -0.029951, -0.047969, -0.037184, -0.004913, 0.032276, 0.032991, 0.009270, 0.018666, -0.031291, 0.002185, -0.007146, -0.054427, -0.034521, 0.027713, 0.037280, 0.030235, 0.007947, -0.057762, -0.179910, -0.126661, -0.035230, 0.107996, 0.016297, 0.016030, -0.025502, -0.028574, -0.017716, -0.045501, -0.035103, 0.014486, -0.031075, 0.015673, -0.009271, -0.012773, 0.019752, -0.000944, -0.044680, 0.015847, -0.031101, 0.036406, 0.028469, 0.114302, 0.140455, 0.139064, 0.076609, -0.093545, -0.173437, -0.044371, 0.108457, 0.123127, 0.090576, -0.001548, -0.059077, -0.062663, -0.019158, -0.049441, 0.003502, -0.041905, -0.000226, -0.024737, 0.012657, 0.028289, 0.010910, -0.018040, -0.043600, -0.022021, 0.003616, 0.098599, 0.091941, 0.171644, 0.241342, 0.198651, 0.034104, -0.079430, -0.127827, 0.004354, 0.125248, 0.146662, 0.094003, 0.005842, -0.018369, -0.042444, -0.008078, -0.020520, -0.016642, 0.004883, -0.029108, 0.001167, 0.016379, -0.033718, -0.020878, 0.018212, 0.000837, 0.020572, 0.083670, 0.119148, 0.202601, 0.215430, 0.245341, 0.226669, 0.044373, -0.043948, -0.059823, 0.013612, 0.171702, 0.148692, 0.087204, 0.021198, 0.052081, 0.015738, -0.036204, -0.000249, -0.009395, 0.031354, 0.019287, -0.021206, 0.031833, -0.006510, -0.008900, 0.010578, 0.051452, 0.066856, 0.096107, 0.180114, 0.251667, 0.226599, 0.229732, 0.168062, 0.086882, -0.001072, 0.004178, 0.096176, 0.232944, 0.243680, 0.151230, 0.130143, 0.094326, 0.002645, 0.025981, -0.027119, 0.020795, -0.018206, 0.006307, -0.000415, 0.016567, 0.005543, -0.025817, 0.016986, 0.040247, 0.049363, 0.118345, 0.174015, 0.208495, 0.208559, 0.195080, 0.167713, 0.109949, 0.089772, 0.089577, 0.157251, 0.246080, 0.217517, 0.157536, 0.094662, 0.080543, 0.005309, 0.022128, 0.021576, -0.037423, -0.024388, -0.028814, 0.009456, 0.006900, -0.018444, 0.021279, 0.013534, -0.026131, 0.046962, 0.098033, 0.155630, 0.201116, 0.151549, 0.098174, 0.134475, 0.074277, 0.097008, 0.177200, 0.273066, 0.293266, 0.195895, 0.149479, 0.049715, 0.031896, -0.005641, -0.005637, -0.040393, -0.005588, 0.010785, 0.025691, -0.006160, 0.032629, -0.033749, -0.010157, 0.005286, -0.000777, 0.026282, 0.023011, 0.101065, 0.054467, 0.040688, 0.036806, 0.004317, 0.033171, 0.088312, 0.207466, 0.221165, 0.178118, 0.105619, 0.018008, -0.039020, -0.057147, -0.076089, -0.023293, -0.044019, -0.028592, -0.039251, 0.004167, -0.005548, -0.024365, 0.022892, 0.029807, -0.035579, -0.003570, -0.032738, -0.027149, -0.006843, -0.033453, -0.022140, -0.059961, -0.088713, -0.022701, 0.029878, 0.117405, 0.090186, 0.052286, -0.018713, -0.080650, -0.102000, -0.046904, -0.053663, -0.030865, -0.053783, -0.032660, -0.019216, 0.000365, -0.025653, 0.005236, -0.022976, 0.005101, 0.024275, -0.021000, -0.022276, -0.102103, -0.108746, -0.153258, -0.159179, -0.180592, -0.156830, -0.113465, -0.023529, 0.022874, 0.017937, -0.031114, -0.012244, -0.045389, -0.109472, -0.081727, -0.045585, -0.088741, -0.060182, 0.006305, -0.005198, 0.011084, -0.014854, 0.006475, 0.023658, -0.009203, -0.019137, -0.059081, -0.057831, -0.067892, -0.165858, -0.172153, -0.165474, -0.200205, -0.164866, -0.113636, -0.086271, -0.048881, -0.069908, -0.016906, -0.048901, -0.063655, -0.072852, -0.043367, -0.070382, -0.066719, -0.043893, -0.033906, -0.020151, 0.027968, -0.027630, -0.020994, -0.029117, -0.018459, -0.006640, -0.038694, -0.039019, -0.066288, -0.123064, -0.130873, -0.155298, -0.122986, -0.127257, -0.070421, -0.067513, -0.063832, -0.029991, -0.056064, -0.042267, -0.005660, -0.013748, 0.005168, -0.025241, -0.022016, 0.015942, -0.003369, 0.031517, -0.018427, -0.011718, 0.001543, 0.019048, -0.031589, -0.013326, 0.015681, -0.018793, -0.026726, -0.092695, -0.125397, -0.138669, -0.125488, -0.114270, -0.062326, -0.067905, -0.089062, 0.006203, 0.006363, 0.035196, 0.009933, 0.043896, -0.015865, 0.031201, -0.022123, 0.011427, -0.014542, 0.022335, -0.029962, -0.006964, -0.009640, -0.021356, -0.017631, -0.011183, -0.001512, 0.010398, -0.034470, -0.008976, -0.073074, -0.079691, -0.061513, -0.058711, -0.047403, -0.027331, -0.028777, -0.032123, 0.008922, 0.040309, 0.021803, 0.051010, 0.060174, 0.031299, 0.000879, -0.003843, -0.017701, -0.004129, 0.031343, -0.018362, 0.005714, -0.026204, -0.009782, 0.001760, -0.029293, 0.003296, -0.043300, -0.035054, -0.002216, 0.000817, -0.039026, -0.058714, -0.075670, -0.061966, -0.056321, 0.006282, -0.032630, 0.024537, 0.022914, 0.000913, 0.033365, 0.020149, -0.002708, -0.026059, -0.011514, 0.011584, 0.030934, -0.012052, -0.014842, -0.034895, 0.021944, 0.034808, 0.023980, -0.022941, 0.017890, -0.027764, -0.010514, -0.018798, -0.081079, -0.062152, -0.067927, -0.102899, -0.045128, -0.046415, -0.043150, -0.067625, -0.068952, -0.056550, -0.012078, -0.022361, 0.022159, 0.027958, 0.001951, -0.029311, 0.014165, 0.031961, -0.008970, -0.018691, -0.008355, 0.005111, -0.026783, 0.018267, 0.011880, -0.021277, -0.027513, -0.038234, 0.000029, -0.015856, -0.031834, -0.046753, -0.039676, -0.008764, -0.029803, -0.051941, -0.012505, -0.032509, -0.012097, -0.028210, -0.002820, 0.001708, -0.021666, 0.022955, 0.032985, -0.029873, 0.010349, -0.024672, -0.007098, 0.017108, -0.000629, 0.010749, -0.011852, 0.033095, -0.018032, 0.005415, 0.001544, 0.022064, 0.000767, 0.018031, 0.003510, 0.018525, -0.003713, 0.008062, 0.032136, -0.013504, -0.015284, 0.025511, 0.013278, -0.033749, 0.012702, -0.035027, -0.019390, 0.013977
--  Sum of weights (converted): FFFFFFFF997B8660
    );

    constant weights_n5 : weight_array := (
     x"009A1E8C", x"80420FA7", x"00F7A6DE", x"0122C0B8", x"00E423CA", x"810CB6E4", x"806A6B55", x"0011CCE0", x"00EDCB3C", x"80311400", x"003D1E32", x"0099FE1C", x"80991D09", x"80B17C4B", x"01211784", x"800689D4", x"00CF051E", x"811D48B8", x"806FAC97", x"00CD4B21", x"801C5337", x"00628BA0", x"80F517CC", x"011CC480", x"80920687", x"800ECB30", x"80BFA21C", x"8081CE63", x"80FAD158", x"81001590", x"803BC567", x"80810CD7", x"00D81E4F", x"80016D28", x"00E35EF2", x"803167B6", x"003D3F7D", x"01180CB8", x"80E31C0C", x"80800B64", x"00F7D7D9", x"8045D81A", x"8051B131", x"0014C353", x"809FAA9F", x"0012BD72", x"807B580F", x"005B8043", x"803F1EAC", x"8062781D", x"806E498D", x"004BFEC9", x"0092D2F3", x"810B7B04", x"80CC0C4C", x"8118C936", x"0088923C", x"00DB6BEE", x"81191AD6", x"004BFCA3", x"003B23DC", x"809D0DEB", x"003EDC11", x"00E0020E", x"011C0590", x"00788C4E", x"80460081", x"80BA4332", x"808DCC65", x"802A9271", x"8050F0F2", x"009BBC8A", x"8134B152", x"8006B9CA", x"80769985", x"00003123", x"01008F50", x"800A6357", x"803D5DC6", x"8067FD78", x"812615A2", x"81097C00", x"007F7A97", x"80B2A9EA", x"00A61B45", x"8052F297", x"00698BF2", x"00D55521", x"002BD47D", x"005E8F15", x"00EFC46D", x"806CE5A5", x"00BD3D16", x"81278448", x"00C511B4", x"80D014F1", x"808D4F24", x"80031B4A", x"8098B68C", x"0061C78B", x"810A1AE6", x"80FE1193", x"00DB4306", x"80DB454C", x"00A38E91", x"0106E71E", x"00C429FE", x"807C3057", x"800CA3C1", x"8106F938", x"809EE252", x"803C8E57", x"80C14D21", x"00A8C6DC", x"0099232F", x"80551C67", x"8037D552", x"00F1120C", x"805BD581", x"007C08A5", x"003CA276", x"8168B16C", x"8225620C", x"80284C0E", x"82428F0C", x"810F622C", x"828A2628", x"80F25CCE", x"8014D26D", x"80229F87", x"0150245A", x"80BB3AFB", x"8017B92E", x"00CDBE22", x"01FE1C40", x"017B0962", x"0145A624", x"00A62586", x"0111C3D2", x"80493410", x"805A51FB", x"80282CF2", x"00722555", x"805E875F", x"003981DC", x"80320C1D", x"80954044", x"801B2189", x"80EB8714", x"8026744A", x"80C68C39", x"817309E6", x"804C2C73", x"80FA0C31", x"8062E8FF", x"80898987", x"80152B7A", x"001E9214", x"0078357F", x"020DDE50", x"037F6A38", x"031BEFBC", x"0344A974", x"03BE1A4C", x"0173E858", x"012D3570", x"80BA9BDA", x"8107A826", x"80AAAF8A", x"80321B9E", x"00613C0D", x"0073C903", x"81299B00", x"810BBD26", x"80C26CE9", x"8154E828", x"80B1E141", x"00C4E7D9", x"0097E301", x"01BEEFE4", x"018B5E96", x"007A179A", x"80223087", x"81184B28", x"80CE1654", x"00BA6D11", x"02569FB4", x"036C3CF0", x"037CEB88", x"053198A8", x"04D4EA80", x"05B8D300", x"03C2B63C", x"0271C168", x"01824304", x"0075023F", x"00139A56", x"806C6C96", x"80F7B8B5", x"810345E2", x"81BD112E", x"804DCBD2", x"81ABDF18", x"80DD8BC8", x"80B60B76", x"00D7CF1E", x"030AA1FC", x"02787640", x"01139A6A", x"00BB7BC2", x"0054EC5E", x"80B9E283", x"821D0604", x"80166725", x"000E6C1D", x"015E04B0", x"0416FBD8", x"03897750", x"05271898", x"079F9028", x"07B3E560", x"02A5AE54", x"002192C1", x"80679A75", x"00E2A2F9", x"00A98067", x"00A889A1", x"0066EAD6", x"813B51D8", x"8059262E", x"81259910", x"80362D14", x"00BC9720", x"02303EA4", x"02A5CDC8", x"0247D1B0", x"023C57BC", x"808A9689", x"80D89083", x"80F05451", x"81717EF0", x"81C7AAF8", x"80E3C8A3", x"010948E8", x"02684034", x"04042F98", x"060231E0", x"07C48E38", x"06DD9EA0", x"039E6A40", x"020C4690", x"80150AA8", x"80739BC3", x"80D8C520", x"010A4366", x"0041A53E", x"817C4CBA", x"81EF7BA4", x"005B66D0", x"00DEAB20", x"01BA1B50", x"018B44B8", x"0396970C", x"02E7C7FC", x"030FC124", x"0027C521", x"81230FE0", x"82A191D0", x"8193651C", x"8186A37E", x"83089184", x"803E8C5C", x"8064CD6B", x"00DF20EC", x"03D6FE80", x"05DA6300", x"06C6CAE8", x"0401E118", x"01D5DD64", x"80EE1040", x"00867611", x"805F8B4A", x"800070F1", x"00876B0A", x"8147D99E", x"00055809", x"803734FC", x"01EB9C4E", x"029641A8", x"043C9370", x"05804518", x"04EB6D28", x"03BC3838", x"04692480", x"00B03E35", x"809A0145", x"8242C0F4", x"84CB5580", x"843F2708", x"840E45B0", x"83D25808", x"81F3873E", x"80E4A672", x"022E72F4", x"038B2DF0", x"017814BE", x"00A42B8E", x"00A3114F", x"00DF6355", x"005FE9E4", x"006CB9ED", x"8069B73A", x"803AB350", x"80E61E2F", x"019AD92A", x"02A59304", x"0280FB30", x"03273FE4", x"0632E4C8", x"05F8A1A0", x"07C14280", x"041C0420", x"0166682C", x"81C59D8C", x"82D6A8B4", x"8643A2D0", x"863F2208", x"873A3BC0", x"85E59B58", x"84D72ED0", x"836950FC", x"81216210", x"806DB942", x"006F2D9C", x"0096688B", x"01042F18", x"806BBC26", x"80E94687", x"80F05B93", x"80A09550", x"00172044", x"000159AE", x"0094EB4E", x"01892552", x"03C09AE8", x"0373F31C", x"079A4728", x"08516F20", x"08436D80", x"059E33C8", x"0103B094", x"80D050B1", x"84409B28", x"85302050", x"86D04928", x"8616DFA8", x"85AEC878", x"856F33C0", x"84D74EC8", x"825C68C0", x"807B68D6", x"00C3773F", x"80266015", x"003223EA", x"80CC4872", x"80DC7AD9", x"80396E00", x"0014AEB1", x"80ACD2C1", x"80D46F9B", x"00EDB84A", x"02155728", x"0237792C", x"05947498", x"06448158", x"08C26490", x"0771E9A0", x"03701504", x"0174EC2E", x"83364D20", x"8485CAA0", x"82DC4ADC", x"8338BE70", x"8359E734", x"83392854", x"8403A038", x"82EBA114", x"81EB7F4C", x"80D20EFA", x"001AD22A", x"0047EDAA", x"00068801", x"0023C42D", x"000493EB", x"00C3E318", x"0099213D", x"8039E003", x"8014DAEF", x"80AF459A", x"0023A590", x"023C50AC", x"030B8A44", x"05D3A2B0", x"0531C5E0", x"033E1E94", x"007AE8BC", x"8160CA1C", x"825FB404", x"848DD010", x"82F53DAC", x"812328C4", x"81FC4A06", x"80CCCBD0", x"81F0BAC4", x"836DE9F0", x"8215EEDC", x"820FC6B4", x"00D5BDCE", x"00847B57", x"006FED14", x"00E10F52", x"00DF38E1", x"011FD292", x"00700D47", x"811B6190", x"803EB670", x"81C224A6", x"82CA4950", x"81CE6DEC", x"01596F00", x"01A05A90", x"01FFDE30", x"006DCAB4", x"8081CEC4", x"84178CF0", x"83D7E92C", x"8385E594", x"82C900E8", x"00153401", x"800E6A56", x"806FA6DA", x"805E1985", x"818294DA", x"814C0BE8", x"818EEA9C", x"80253710", x"80907212", x"00A86CF4", x"00FE6DE6", x"811142BC", x"80AE15E4", x"01129D8E", x"80D4DAE7", x"806E32FB", x"813D26B6", x"83C5A7E4", x"85147388", x"83542C0C", x"83037344", x"826CB9E4", x"82F01BBC", x"82B77FB8", x"846FDDE0", x"8327FC48", x"82964D5C", x"810B334A", x"8100060E", x"002D179E", x"806BF153", x"813E805C", x"80206364", x"80565137", x"00349DFD", x"802AB310", x"801134E8", x"800CD6C6", x"009E093E", x"80CAC223", x"0037B896", x"00925A15", x"0069DFB7", x"81048782", x"00914609", x"82E21E1C", x"83B41048", x"84911558", x"85F05490", x"85121C98", x"85DFD888", x"845ABF60", x"835CA338", x"831BCE2C", x"81439CD0", x"006AABC6", x"0053F2B3", x"01CB234A", x"80358D52", x"00C1857C", x"00CC08EA", x"012522C2", x"8055F9E3", x"8129B6D4", x"80722A83", x"00D84BF2", x"00197E6F", x"01175868", x"80DF7BE0", x"80D73716", x"00764139", x"00D00838", x"0180B816", x"01F84A0E", x"823F80F0", x"84CC8060", x"84B2AFE0", x"85495978", x"840DFF10", x"82D0D4C4", x"80D1EF92", x"800B88A8", x"00A246D8", x"80210CD3", x"0069CD86", x"01EAAD56", x"00720AFA", x"002BC84A", x"002E4D9F", x"809059BA", x"8087500E", x"00ECAB35", x"00326D0B", x"0035DBD7", x"0073FBD8", x"00B138C6", x"00BE59E4", x"00983281", x"003E8C03", x"01B163CA", x"043FF1D8", x"035C6DD4", x"0230B0F8", x"80B49EF6", x"824FEEA0", x"8045DE5F", x"816A94EC", x"80B371BA", x"81120964", x"811C8400", x"80002EBF", x"0111F3A8", x"0028E0EA", x"0112F2D6", x"003DEA41", x"010D2140", x"01762A90", x"00465945", x"802FEDB3", x"00B008F2", x"80C0208D", x"803C282F", x"80F39768", x"00CC575E", x"0055B291", x"80BAC008", x"0054848E", x"018160B0", x"038E8F10", x"03B51A08", x"047C3778", x"04935668", x"033860AC", x"015F091E", x"01BE2D70", x"804A749D", x"80419461", x"80006388", x"0015D104", x"004D0E67", x"01F211D6", x"02063F00", x"01F54936", x"00485859", x"00FDC356", x"00AE367D", x"800BCEF1", x"80429F4D", x"806B71CD", x"0064D469", x"008B0764", x"80394000", x"00D9680F", x"803B0FBA", x"8020621B", x"80064E74", x"0106AE84", x"036D1E30", x"0490B810", x"05204588", x"035F7384", x"0279378C", x"00652EB3", x"802EF4A1", x"800D3B08", x"00D8C57A", x"8011889F", x"019B86D0", x"02A05418", x"01031650", x"02469E4C", x"017C3ACE", x"800D82D1", x"00A1FF47", x"80A3429D", x"003D2F31", x"81065C4A", x"0112EA52", x"807CD4E5", x"00BB17A9", x"80C17545", x"811EB6E6", x"00367B07", x"002A1F94", x"80252F36", x"004EE144", x"025E3CF4", x"02C3DAE8", x"03D23704", x"034045BC", x"03212000", x"02FF758C", x"0115DE18", x"02D3A590", x"036B2788", x"02A1F0C8", x"0125164A", x"0104AEE0", x"01B9FE20", x"019CB6D2", x"0108E69E", x"004E6289", x"80A4832B", x"80F808D1", x"80A4EF4A", x"00022CBB", x"00269069", x"00E012C1", x"80D5DE57", x"0089D661", x"00E00958", x"8137B3C4", x"80D2EEB2", x"800BB763", x"01673BBA", x"0306E1E8", x"02DDDD8C", x"03D22168", x"0400BEC0", x"03B5C93C", x"01C526D6", x"01CBBCA2", x"0226B060", x"0174F214", x"00F6E231", x"01953DD0", x"0169B04A", x"80431C1C", x"807D787B", x"002B4680", x"0032044E", x"00BB735B", x"00693FA4", x"005B2B2B", x"00600C82", x"00D9D3F5", x"00AD95D9", x"801F501D", x"80E0F84A", x"009D2B97", x"803B6687", x"80B8BB9B", x"0027194A", x"01DD4534", x"00E1F035", x"01D1CBD8", x"02B0CD50", x"03183AD0", x"01C1AB72", x"00589CDC", x"801E7A01", x"80380430", x"002C59CA", x"80D99B81", x"00E52D79", x"00388848", x"80CB249F", x"00AADFC1", x"001858D8", x"011CC924", x"8005ECA6", x"8003DBB9", x"811A5E04", x"80F1A941", x"0001023B", x"00FAD711", x"80B68706", x"0021D9EA", x"80F111E5", x"81063BA0", x"808CBE38", x"80B7A3B4", x"80CD7035", x"8007BC7D", x"00309DDB", x"00CE5C03", x"0063C13E", x"8040176E", x"808C1A70", x"807ACA12", x"8132D2F0", x"00904DF9", x"00D82700", x"81117626", x"8105F156", x"81010F22", x"8024807F", x"8000C635", x"80BF0C0E", x"00A1AB13", x"0013447D", x"8094175E", x"811B08C0", x"00E3C260", x"011F10C0", x"0013921C", x"809BE640", x"009BDA47", x"007D0C8C", x"8060BF09", x"00D51D3B", x"81153B30", x"80617C63", x"00A19290", x"8117F4CE", x"80A092AB", x"80C12D0E", x"80B63954", x"00C79CB7", x"009111BF", x"8116B548", x"80B442DD", x"80026E11", x"805F931D", x"80A1381D", x"811F9E68", x"00D7C75A", x"00A3CE90", x"0054E42B", x"8041D790", x"811B987C", x"80125104", x"006FD712", x"80553E97", x"00E58278", x"00415E7C", x"801103F9", x"00707174", x"009627A6", x"80D72176", x"0053A3CA", x"8116E5C8", x"804F615A", x"806D1423", x"00D1709D", x"812759CC", x"005D2299", x"8110B820", x"007C2F8A", x"004680A3", x"8074098A", x"005651E8", x"0118CD36", x"00B21EA3", x"810AF644", x"804BD272"
--  0.018813, -0.008064, 0.030231, 0.035492, 0.027849, -0.032802, -0.012991, 0.002173, 0.029028, -0.005991, 0.007461, 0.018798, -0.018691, -0.021666, 0.035290, -0.000798, 0.025271, -0.034825, -0.013632, 0.025060, -0.003458, 0.012029, -0.029919, 0.034762, -0.017825, -0.001806, -0.023393, -0.015845, -0.030617, -0.031260, -0.007296, -0.015753, 0.026382, -0.000174, 0.027755, -0.006031, 0.007477, 0.034186, -0.027723, -0.015630, 0.030254, -0.008526, -0.009972, 0.002535, -0.019491, 0.002288, -0.015057, 0.011170, -0.007705, -0.012020, -0.013463, 0.009277, 0.017923, -0.032651, -0.024908, -0.034276, 0.016671, 0.026785, -0.034315, 0.009276, 0.007219, -0.019172, 0.007673, 0.027345, 0.034671, 0.014715, -0.008545, -0.022737, -0.017309, -0.005197, -0.009881, 0.019011, -0.037682, -0.000821, -0.014478, 0.000023, 0.031318, -0.001268, -0.007491, -0.012694, -0.035899, -0.032408, 0.015561, -0.021810, 0.020277, -0.010125, 0.012884, 0.026042, 0.005350, 0.011543, 0.029268, -0.013293, 0.023100, -0.036074, 0.024056, -0.025401, -0.017250, -0.000379, -0.018642, 0.011936, -0.032484, -0.031014, 0.026765, -0.026766, 0.019965, 0.032093, 0.023946, -0.015160, -0.001543, -0.032101, -0.019395, -0.007392, -0.023596, 0.020603, 0.018694, -0.010390, -0.006816, 0.029428, -0.011210, 0.015141, 0.007402, -0.044030, -0.067063, -0.004919, -0.070625, -0.033128, -0.079364, -0.029585, -0.002542, -0.004226, 0.041033, -0.022855, -0.002896, 0.025115, 0.062269, 0.046269, 0.039752, 0.020282, 0.033419, -0.008936, -0.011025, -0.004904, 0.013934, -0.011539, 0.007020, -0.006109, -0.018219, -0.003312, -0.028751, -0.004694, -0.024237, -0.045293, -0.009299, -0.030523, -0.012074, -0.016789, -0.002584, 0.003732, 0.014674, 0.064193, 0.109304, 0.097160, 0.102132, 0.116956, 0.045399, 0.036769, -0.022779, -0.032185, -0.020836, -0.006117, 0.011869, 0.014134, -0.036329, -0.032683, -0.023734, -0.041615, -0.021714, 0.024036, 0.018541, 0.054558, 0.048263, 0.014904, -0.004174, -0.034216, -0.025157, 0.022757, 0.073074, 0.106963, 0.108999, 0.162304, 0.150991, 0.178812, 0.117519, 0.076386, 0.047151, 0.014283, 0.002393, -0.013235, -0.030239, -0.031650, -0.054329, -0.009497, -0.052230, -0.027044, -0.022222, 0.026344, 0.095048, 0.077205, 0.033643, 0.022886, 0.010367, -0.022691, -0.066043, -0.002735, 0.001761, 0.042727, 0.127806, 0.110531, 0.161022, 0.238228, 0.240710, 0.082725, 0.004098, -0.012647, 0.027666, 0.020691, 0.020573, 0.012563, -0.038491, -0.010882, -0.035840, -0.006613, 0.023021, 0.068389, 0.082740, 0.071267, 0.069866, -0.016917, -0.026436, -0.029337, -0.045104, -0.055624, -0.027806, 0.032383, 0.075226, 0.125511, 0.187768, 0.242744, 0.214553, 0.113088, 0.063998, -0.002569, -0.014112, -0.026461, 0.032503, 0.008013, -0.046423, -0.060484, 0.011157, 0.027181, 0.053968, 0.048251, 0.112133, 0.090794, 0.095673, 0.004855, -0.035530, -0.082223, -0.049243, -0.047685, -0.094796, -0.007635, -0.012305, 0.027237, 0.119994, 0.182909, 0.211767, 0.125229, 0.057357, -0.029060, 0.016414, -0.011663, -0.000054, 0.016531, -0.040021, 0.000652, -0.006739, 0.060011, 0.080842, 0.132395, 0.171908, 0.153739, 0.116726, 0.137835, 0.021514, -0.018799, -0.070649, -0.149821, -0.132709, -0.126742, -0.119427, -0.060978, -0.027911, 0.068170, 0.110740, 0.045908, 0.020040, 0.019906, 0.027269, 0.011708, 0.013272, -0.012905, -0.007166, -0.028091, 0.050152, 0.082712, 0.078245, 0.098541, 0.193713, 0.186601, 0.242341, 0.128420, 0.043751, -0.055373, -0.088703, -0.195756, -0.195207, -0.225859, -0.184278, -0.151267, -0.106606, -0.035325, -0.013394, 0.013572, 0.018360, 0.031761, -0.013151, -0.028476, -0.029341, -0.019602, 0.002823, 0.000165, 0.018179, 0.047991, 0.117261, 0.107904, 0.237583, 0.259941, 0.258231, 0.175562, 0.031700, -0.025429, -0.132886, -0.162125, -0.212926, -0.190292, -0.177586, -0.169824, -0.151283, -0.073780, -0.015065, 0.023861, -0.004684, 0.006121, -0.024937, -0.026914, -0.007010, 0.002525, -0.021097, -0.025932, 0.029019, 0.065105, 0.069272, 0.174372, 0.195862, 0.273730, 0.232655, 0.107432, 0.045523, -0.100379, -0.141332, -0.089391, -0.100677, -0.104725, -0.100727, -0.125443, -0.091263, -0.059997, -0.025642, 0.003274, 0.008780, 0.000797, 0.004366, 0.000559, 0.023912, 0.018693, -0.007065, -0.002546, -0.021395, 0.004351, 0.069863, 0.095159, 0.182084, 0.162326, 0.101333, 0.015004, -0.043065, -0.074183, -0.142311, -0.092437, -0.035542, -0.062047, -0.025000, -0.060636, -0.107167, -0.065177, -0.064426, 0.026091, 0.016172, 0.013663, 0.027473, 0.027249, 0.035135, 0.013678, -0.034592, -0.007655, -0.054949, -0.087193, -0.056449, 0.042167, 0.050824, 0.062484, 0.013402, -0.015846, -0.127875, -0.120106, -0.110095, -0.087037, 0.002588, -0.001760, -0.013629, -0.011487, -0.047190, -0.040533, -0.048696, -0.004543, -0.017633, 0.020560, 0.031058, -0.033357, -0.021251, 0.033522, -0.025983, -0.013452, -0.038715, -0.117878, -0.158746, -0.104025, -0.094171, -0.075772, -0.091810, -0.084900, -0.138656, -0.098631, -0.080847, -0.032617, -0.031253, 0.005504, -0.013177, -0.038880, -0.003954, -0.010537, 0.006423, -0.005212, -0.002100, -0.001567, 0.019292, -0.024751, 0.006802, 0.017865, 0.012924, -0.031803, 0.017734, -0.090102, -0.115730, -0.142710, -0.185587, -0.158461, -0.183575, -0.136078, -0.105058, -0.097144, -0.039503, 0.013021, 0.010248, 0.056047, -0.006537, 0.023623, 0.024907, 0.035783, -0.010495, -0.036342, -0.013936, 0.026403, 0.003112, 0.034100, -0.027281, -0.026271, 0.014435, 0.025395, 0.046963, 0.061559, -0.070252, -0.149964, -0.146812, -0.165204, -0.126709, -0.087992, -0.025627, -0.001408, 0.019809, -0.004034, 0.012915, 0.059897, 0.013921, 0.005345, 0.005652, -0.017621, -0.016518, 0.028890, 0.006156, 0.006575, 0.014158, 0.021634, 0.023236, 0.018579, 0.007635, 0.052904, 0.132806, 0.105033, 0.068444, -0.022048, -0.072257, -0.008529, -0.044260, -0.021905, -0.033452, -0.034731, -0.000022, 0.033441, 0.004990, 0.033563, 0.007558, 0.032853, 0.045675, 0.008587, -0.005851, 0.021489, -0.023453, -0.007343, -0.029735, 0.024944, 0.010461, -0.022797, 0.010317, 0.047043, 0.111152, 0.115857, 0.140163, 0.142986, 0.100632, 0.042851, 0.054465, -0.009089, -0.008005, -0.000047, 0.002663, 0.009406, 0.060800, 0.063262, 0.061192, 0.008831, 0.030977, 0.021266, -0.001441, -0.008133, -0.013116, 0.012308, 0.016971, -0.006989, 0.026539, -0.007210, -0.003953, -0.000770, 0.032066, 0.107070, 0.142666, 0.160189, 0.105402, 0.077297, 0.012351, -0.005732, -0.001615, 0.026461, -0.002140, 0.050235, 0.082071, 0.031627, 0.071120, 0.046415, -0.001649, 0.019775, -0.019929, 0.007469, -0.032026, 0.033559, -0.015238, 0.022838, -0.023615, -0.034999, 0.006650, 0.005142, -0.004539, 0.009629, 0.074004, 0.086408, 0.119411, 0.101596, 0.097794, 0.093684, 0.033919, 0.088336, 0.106830, 0.082268, 0.035777, 0.031822, 0.053954, 0.050380, 0.032337, 0.009568, -0.020082, -0.030278, -0.020134, 0.000265, 0.004708, 0.027353, -0.026107, 0.016826, 0.027348, -0.038050, -0.025749, -0.001430, 0.043852, 0.094590, 0.089583, 0.119401, 0.125091, 0.115941, 0.055316, 0.056120, 0.067223, 0.045526, 0.030137, 0.049468, 0.044151, -0.008192, -0.015316, 0.005283, 0.006106, 0.022882, 0.012848, 0.011129, 0.011725, 0.026590, 0.021190, -0.003822, -0.027462, 0.019186, -0.007251, -0.022550, 0.004773, 0.058261, 0.027580, 0.056860, 0.084082, 0.096708, 0.054891, 0.010817, -0.003720, -0.006838, 0.005414, -0.026563, 0.027976, 0.006901, -0.024798, 0.020859, 0.002972, 0.034764, -0.000723, -0.000471, -0.034469, -0.029500, 0.000123, 0.030620, -0.022281, 0.004132, -0.029427, -0.032011, -0.017181, -0.022417, -0.025078, -0.000944, 0.005935, 0.025190, 0.012177, -0.007824, -0.017102, -0.014989, -0.037454, 0.017615, 0.026386, -0.033382, -0.031975, -0.031379, -0.004456, -0.000095, -0.023321, 0.019735, 0.002352, -0.018078, -0.034550, 0.027803, 0.035042, 0.002389, -0.019031, 0.019025, 0.015265, -0.011810, 0.026015, -0.033842, -0.011900, 0.019723, -0.034174, -0.019601, -0.023581, -0.022244, 0.024367, 0.017709, -0.034022, -0.022005, -0.000297, -0.011667, -0.019680, -0.035110, 0.026340, 0.019996, 0.010363, -0.008037, -0.034619, -0.002236, 0.013652, -0.010406, 0.028016, 0.007980, -0.002077, 0.013726, 0.018329, -0.026261, 0.010210, -0.034045, -0.009690, -0.013315, 0.025566, -0.036054, 0.011369, -0.033291, 0.015159, 0.008606, -0.014165, 0.010537, 0.034278, 0.021743, -0.032588, -0.009256
--  Sum of weights (converted): 000000009FD127B4
    );

    constant weights_n6 : weight_array := (
     x"01096320", x"002D43AB", x"002411CD", x"0014DFCD", x"8066DD25", x"804C88B7", x"00136AB2", x"00DC3BE3", x"805275F5", x"804C905E", x"0037B19E", x"806B1530", x"01007DA8", x"00DE78C7", x"000BCA99", x"80BD37D6", x"0051E18B", x"00F81D95", x"00606282", x"007AA225", x"809ADCB5", x"812036D4", x"806E03D5", x"00095999", x"0103F0EE", x"003D1660", x"8035A25D", x"80498419", x"8037F0DB", x"809D52FE", x"807A7C3E", x"00365A84", x"00C636D9", x"00F8C8E5", x"0076549A", x"80BB4E40", x"0123F206", x"013724D6", x"802D9193", x"00425CE7", x"014C4380", x"80344235", x"00AB187E", x"004ECCF3", x"00BF4EFC", x"0085571A", x"013BE842", x"010AA406", x"80B8BA32", x"00B8BA88", x"803571E8", x"80979DEF", x"0031124D", x"8027D299", x"80BEA91A", x"81023F2E", x"80A30DA7", x"001E1F3D", x"00B2507C", x"00AC61F3", x"005187D3", x"0116C828", x"80EDA2E3", x"808AA62E", x"00D0A7DC", x"807C154F", x"020CDFC0", x"016EF97A", x"013220B8", x"02DCB428", x"028486F4", x"02DC936C", x"02BBDBA4", x"01A3C7A8", x"02BBAFEC", x"01927704", x"0114087C", x"010BCBC2", x"8080E770", x"80882CCB", x"011E50CA", x"80BF4636", x"009E1643", x"00B0D237", x"80ED8631", x"802187E9", x"80032875", x"00D9C072", x"804CFDA7", x"010BF06E", x"80DA9C42", x"00BBE9D9", x"011C1870", x"0069ADAA", x"00F48AB8", x"00FA0562", x"025413F4", x"02F77BE4", x"02EABED0", x"04D9C000", x"045187E0", x"04D4EC38", x"05CC29F0", x"04B54FD8", x"03FD958C", x"02F7C2F0", x"008BB2E9", x"00A22C49", x"014D2946", x"80ABF3F0", x"0028CB73", x"00D9547C", x"00204DC7", x"80419A8E", x"00699DE9", x"80F263A6", x"00F0D08F", x"00DE36B7", x"8056F44A", x"8061BFD9", x"000A4819", x"019D20F0", x"004531D6", x"00C7CC4C", x"809E7207", x"0128F964", x"01F6777E", x"026553D4", x"0345C554", x"04AE84B0", x"060D86E8", x"05471940", x"037847E0", x"01B21894", x"025D5AA4", x"00540FD7", x"00FC16B7", x"802D3812", x"0003FDF9", x"80E54368", x"806F7579", x"001823CB", x"811A93B6", x"80416FD1", x"00A0D9C2", x"009D6971", x"0085E4E6", x"80BBF1F8", x"800B20F2", x"810BD170", x"004F7AA5", x"80CE6A9A", x"801CCBE1", x"817FDC54", x"0001561A", x"0019D748", x"0193942A", x"019CB21E", x"015D32A4", x"013F0C2E", x"00531EFF", x"00F93628", x"8090A33D", x"80428367", x"009A739F", x"0105A0B6", x"804A3B4D", x"00CCA09D", x"80162B84", x"803A8CA1", x"80233D5F", x"8093B8F3", x"002BA73E", x"805AA1FF", x"812A83D0", x"001F6820", x"811F037A", x"8179AA44", x"80D81880", x"81B8B1E8", x"8278DA24", x"836C17A4", x"82F88E94", x"82F19288", x"81206F1A", x"81EDA552", x"815F30C0", x"816D52FC", x"81E0C630", x"81E75E10", x"81E88B1E", x"80B5E4C4", x"818FAB46", x"80CAC0C4", x"00DA5072", x"8037E65F", x"00EC062C", x"00AD2C72", x"803F3A84", x"81044DEA", x"00ADFC9E", x"8071DA94", x"003324A4", x"81D271D8", x"80A728D5", x"81FFB108", x"81CD1838", x"83023C88", x"8392577C", x"831F28FC", x"81D77D50", x"829BB528", x"83D915F8", x"83CA58CC", x"8587E6F8", x"86148C60", x"83EDC540", x"82E1F210", x"81C08EA4", x"80F91E05", x"00148E90", x"80E2C538", x"00103B40", x"806AE0A2", x"8026F71A", x"00E715E4", x"80EC2F2D", x"007F483E", x"80FE3CF6", x"80BE2659", x"8133610E", x"816A6BE2", x"80C574C7", x"819F96EE", x"80C51119", x"82609C04", x"81CED708", x"82CB3368", x"831713E4", x"82622E38", x"859EFCB0", x"87A13CA0", x"87F4F508", x"8754A028", x"859FC2C0", x"84F0B2C0", x"83C2466C", x"81A3424A", x"80CBD87A", x"00688D73", x"80037155", x"804E81C7", x"803E9EFD", x"803C5560", x"806433CE", x"808F8708", x"80BBF262", x"807B267D", x"807F566D", x"003BF1D1", x"8180964E", x"80188641", x"8178E296", x"8299AB84", x"809509BC", x"817701C6", x"81A904FE", x"836C5C60", x"865C8600", x"8789F3D8", x"89315740", x"86BA8E28", x"8538B5C0", x"83AA04E4", x"8385D4EC", x"81BA342A", x"80D356B3", x"007CCFEA", x"80D748C2", x"810FA48C", x"81090624", x"00258762", x"80E81F61", x"80621C09", x"80F880F4", x"80855C08", x"816DA5FA", x"009B537F", x"8101779E", x"8108709C", x"80407810", x"8197931C", x"007D153A", x"00633CCC", x"81F8550E", x"8404E6C8", x"874CF550", x"870FBE88", x"87317F78", x"8549CD68", x"83470A14", x"81A7A300", x"82476AC4", x"81F48DF0", x"8165CE9E", x"8018EA2D", x"0055F309", x"0095CA75", x"007EE4A7", x"011ACBCA", x"80E46026", x"810E7984", x"80C207CB", x"006A2B67", x"810C0696", x"01494690", x"00BD1811", x"0127F850", x"0158BDCA", x"01C58252", x"02EE9F50", x"00D497DD", x"8306CDD4", x"84FC06A0", x"8467BDB0", x"84C304F8", x"84595AF8", x"835920F0", x"82295ABC", x"0076ABF2", x"80567832", x"01E0A918", x"00266CD4", x"80DACEBE", x"8080C07D", x"80B51979", x"80FE4077", x"001C5501", x"804702E5", x"80A60D0D", x"809D38FC", x"80858F56", x"00BE1F2B", x"8016610D", x"00FD53C5", x"00EB3C62", x"00123807", x"0337F73C", x"02052BFC", x"00F2A2AB", x"8294D77C", x"83EF68DC", x"81BF4FE0", x"82E9D768", x"81E20330", x"81FA57E8", x"803A0706", x"02552724", x"03703614", x"01ACDC64", x"00A82FF9", x"809DD0D1", x"802F2416", x"80F47D22", x"80E793C6", x"8040ACD8", x"0116BC9E", x"0016656A", x"80E67567", x"008376F8", x"015528C4", x"01CCF998", x"0170DFC4", x"01783112", x"03105AFC", x"03BD63D4", x"02D577B4", x"804ED679", x"82AD2794", x"000AC943", x"0066EB16", x"010779F2", x"009C9DE4", x"012B6490", x"0242A694", x"03EB1E38", x"031A4E04", x"02DD6AE8", x"01809794", x"80775563", x"00BD039D", x"0016D36F", x"804A2A72", x"80835627", x"81057F72", x"8001BB32", x"007D1088", x"006764A1", x"016772CA", x"021933C4", x"02493BB8", x"0286B008", x"029E59B4", x"047B4420", x"00750291", x"81DD80EC", x"0025F682", x"023FBF18", x"018FB93A", x"01437D6A", x"816A48F8", x"00B29F00", x"027EE8D0", x"03A976B4", x"035A4B08", x"028E0E78", x"02A796AC", x"006F76DD", x"80A22DF8", x"01191A80", x"803D17F6", x"8036246F", x"004A2017", x"00D01169", x"8129BF22", x"809780B3", x"801BB255", x"00EEA0D6", x"02101D50", x"03853098", x"05385288", x"031EEBF4", x"01CDE6EC", x"00F52484", x"0189F790", x"0237E898", x"01A3C42A", x"81116D5A", x"00688B86", x"0057771D", x"024631E0", x"042AEB10", x"041716F8", x"022807C0", x"0079D7CD", x"80FC416F", x"8126C960", x"80414312", x"80E3261F", x"801D9BA8", x"809DF3CC", x"0074C97A", x"8002F214", x"0009A357", x"80CB7877", x"00B225B8", x"032F75A8", x"045124D0", x"069CE9D8", x"03C31D8C", x"02B676B4", x"0041DE41", x"009699DD", x"00786836", x"816EEE36", x"8201A658", x"00B1F9B2", x"02477220", x"032BFFE0", x"03248980", x"02ACCFE0", x"011C0A2C", x"01BBC582", x"80C64E2F", x"81336CFA", x"00F24B42", x"80179870", x"00C477C2", x"806658EC", x"00A263F2", x"81CF084A", x"80BC1CD5", x"000E1BF8", x"0133C7E2", x"04082C88", x"0565CFD8", x"060F5BE8", x"06901898", x"022FBC70", x"0182CEA2", x"808BF3B9", x"81AFEA9E", x"82108594", x"80BF73B5", x"00B5CD81", x"02722FB8", x"020F3C84", x"01DC083A", x"00DA45D9", x"0020E07A", x"8066B189", x"00ADA02A", x"80F72047", x"80E26065", x"80EE32DD", x"01119D78", x"802AED02", x"80A13E24", x"80803FFD", x"829321C0", x"81ED6538", x"0166AA42", x"0394F564", x"04CFAA88", x"07A337A8", x"0789F740", x"0557A7F8", x"0194590C", x"011AD228", x"8020F9A0", x"80210CB0", x"02F160B0", x"02E7A7F0", x"03C9926C", x"01E1433E", x"01E2CA68", x"009E230E", x"81221154", x"80F2BBDE", x"80513F70", x"80BDA204", x"00241AC0", x"009A7EE4", x"00220096", x"81271426", x"8058F5F8", x"81A9DB76", x"81C1CDF6", x"83114178", x"81B0EC8E", x"01521BEE", x"05082678", x"074998C8", x"086E4C90", x"06AC2190", x"0309FA50", x"026F06C8", x"02F3210C", x"044C2450", x"053BE3C8", x"04ACC4F0", x"03D95260", x"01E925E2", x"0058ED61", x"00AC64C5", x"001A8727", x"80163FED", x"00771922", x"0075298A", x"00FF4F39", x"00FE81EA", x"80EEAD01", x"811B9570", x"80E4009C", x"802820AC", x"80FCA61D", x"8294F8CC", x"8301FB48", x"816081EE", x"0248B4BC", x"0646C948", x"07BE9298", x"07376D98", x"080C2B40", x"075E2390", x"059A8080", x"0501ACA8", x"050EDFA0", x"024DE6B4", x"026A2644", x"8002B013", x"80D4A41E", x"81C3A2C4", x"82093DA4", x"804C8FA7", x"809B5C66", x"80B4585C", x"00E9354C", x"00364047", x"804E82B5", x"81133BB0", x"80D3CADB", x"81165958", x"81258E2A", x"83A2C114", x"824A4C20", x"818D82FE", x"810829F4", x"8015FCE1", x"03E71F48", x"05608A78", x"06DECEC8", x"05EE4708", x"0528D9D8", x"02D34D10", x"01AF52FE", x"00A2F754", x"81BFE054", x"813A4774", x"8069A544", x"8038E16C", x"808A579B", x"80826B1A", x"005EA890", x"81044A24", x"80581EE8", x"00FDC3FC", x"0025A647", x"8006541A", x"80FC9E70", x"811858B6", x"80C7E020", x"82B62500", x"831AD654", x"841BC238", x"83A4CB1C", x"8373C134", x"840E0270", x"8182EE54", x"8177FB8E", x"821B00E4", x"8104E6AC", x"830AE024", x"838DD440", x"825E41C0", x"82B92E08", x"820D3E54", x"8216C5F8", x"81026BEE", x"00817D46", x"8132B4FE", x"80D16916", x"8040F796", x"80E78C33", x"0036C3F2", x"803A23B0", x"00DCABE1", x"812A9010", x"80166FF3", x"00238D64", x"80AC46F9", x"81E64522", x"8184073E", x"84869608", x"83B840EC", x"854D1060", x"856AF160", x"8502BB90", x"855F0230", x"84B6D818", x"844742E0", x"84414468", x"81C28EF0", x"80A83D01", x"808E405E", x"80D562E4", x"8162AAA8", x"80366AC7", x"00373164", x"80E9F35F", x"00F845BF", x"8007B454", x"004FE892", x"01021A26", x"007EF608", x"809F7D58", x"00640C00", x"008FD70C", x"004B4037", x"811BC188", x"80E842F0", x"826109AC", x"82448C1C", x"837672B8", x"8249DC04", x"81E96AEC", x"83F6E648", x"830073A4", x"827C2754", x"825DE0FC", x"801D6851", x"81B1C8E4", x"8120513A", x"81443F02", x"802CFA9D", x"80ED8C7C", x"80CB73D8", x"01221B02", x"0082ABB0", x"007C1F29", x"00CF7D9A", x"00328DA9", x"002F7896", x"80DBEB33", x"00502C13", x"80ECDD3F", x"8017EC85", x"80CD29B2", x"80F97698", x"81287940", x"813C7394", x"817A9380", x"817E3D76", x"81517CF0", x"81ED4E48", x"001D7ACE", x"8053214E", x"81B9E760", x"819632FC", x"80E0E0DD", x"003FA8DC", x"00EE6DF9", x"803C363B", x"00A652F5", x"80A04DED", x"803CC700", x"802D6488", x"811CD826", x"000186C0", x"004D6F0E", x"00B25345", x"80E27110", x"8058EF7B", x"0009471D", x"0019403F", x"00256FEE", x"80EE7F6D", x"00C5BC7A", x"813358CA", x"809AE2C4", x"005778E1", x"80864F1D", x"80C704E6", x"8153E9F6", x"00981435", x"80343C3E", x"006AE687", x"00160792", x"80EABF5A", x"80706A62", x"00CDF76E", x"808FC407", x"8086E557", x"00A06C75", x"807ECCE2", x"002FC2B4", x"808E3B85", x"005A0EF0", x"001DC302", x"80E83B1A", x"80DDE8F5", x"006B69D9", x"80604805", x"009F8F4B", x"000E17E7", x"80658E39", x"803528AB", x"8087E98F", x"008BA808", x"00E1C62B", x"80110A5E", x"80C2EEE0", x"00CBC8A7", x"00E752B8", x"00C2B54A", x"80082A95", x"004652D6", x"000DE6C5", x"80701B40", x"8121C410", x"8023C2B7", x"007E89C9", x"00AAA91C", x"004595C2"
--  0.032396, 0.005525, 0.004403, 0.002548, -0.012557, -0.009343, 0.002370, 0.026884, -0.010066, -0.009346, 0.006799, -0.013072, 0.031310, 0.027157, 0.001439, -0.023098, 0.009995, 0.030288, 0.011766, 0.014970, -0.018904, -0.035182, -0.013430, 0.001141, 0.031731, 0.007457, -0.006547, -0.008974, -0.006829, -0.019205, -0.014952, 0.006635, 0.024196, 0.030369, 0.014445, -0.022864, 0.035638, 0.037981, -0.005563, 0.008101, 0.040560, -0.006379, 0.020886, 0.009619, 0.023353, 0.016277, 0.038563, 0.032549, -0.022550, 0.022550, -0.006524, -0.018508, 0.005990, -0.004861, -0.023274, -0.031524, -0.019904, 0.003677, 0.021767, 0.021043, 0.009952, 0.034031, -0.029008, -0.016925, 0.025471, -0.015147, 0.064072, 0.044797, 0.037369, 0.089441, 0.078678, 0.089426, 0.085432, 0.051243, 0.085411, 0.049129, 0.033695, 0.032690, -0.015735, -0.016623, 0.034951, -0.023349, 0.019298, 0.021585, -0.028995, -0.004093, -0.000386, 0.026581, -0.009398, 0.032707, -0.026686, 0.022939, 0.034680, 0.012900, 0.029851, 0.030520, 0.072763, 0.092710, 0.091155, 0.151581, 0.134952, 0.150992, 0.181172, 0.147133, 0.124705, 0.092744, 0.017053, 0.019797, 0.040669, -0.020990, 0.004980, 0.026530, 0.003943, -0.008008, 0.012893, -0.029589, 0.029396, 0.027126, -0.010615, -0.011932, 0.001255, 0.050431, 0.008447, 0.024389, -0.019341, 0.036252, 0.061336, 0.074869, 0.102267, 0.146304, 0.189151, 0.164929, 0.108433, 0.052990, 0.073896, 0.010261, 0.030773, -0.005520, 0.000487, -0.027986, -0.013606, 0.002947, -0.034494, -0.007988, 0.019635, 0.019215, 0.016344, -0.022943, -0.001358, -0.032693, 0.009702, -0.025197, -0.003515, -0.046858, 0.000163, 0.003154, 0.049265, 0.050378, 0.042627, 0.038946, 0.010147, 0.030421, -0.017656, -0.008119, 0.018854, 0.031937, -0.009061, 0.024979, -0.002706, -0.007147, -0.004302, -0.018033, 0.005329, -0.011064, -0.036440, 0.003834, -0.035036, -0.046102, -0.026379, -0.053796, -0.077252, -0.106945, -0.092841, -0.091989, -0.035209, -0.060259, -0.042870, -0.044595, -0.058688, -0.059493, -0.059637, -0.022204, -0.048788, -0.024750, 0.026650, -0.006824, 0.028812, 0.021139, -0.007718, -0.031775, 0.021239, -0.013898, 0.006243, -0.056939, -0.020405, -0.062462, -0.056286, -0.094023, -0.111614, -0.097554, -0.057555, -0.081507, -0.120250, -0.118451, -0.172840, -0.190008, -0.122775, -0.090081, -0.054756, -0.030410, 0.002509, -0.027682, 0.001981, -0.013047, -0.004757, 0.028209, -0.028831, 0.015537, -0.031035, -0.023212, -0.037522, -0.044241, -0.024104, -0.050731, -0.024056, -0.074293, -0.056499, -0.087305, -0.096567, -0.074485, -0.175658, -0.238432, -0.248652, -0.229080, -0.175752, -0.154382, -0.117465, -0.051179, -0.024883, 0.012763, -0.000420, -0.009583, -0.007644, -0.007365, -0.012232, -0.017520, -0.022943, -0.015033, -0.015544, 0.007317, -0.046947, -0.002994, -0.046006, -0.081259, -0.018193, -0.045777, -0.051882, -0.106978, -0.198794, -0.235590, -0.287273, -0.210273, -0.163173, -0.114504, -0.110087, -0.053980, -0.025798, 0.015236, -0.026280, -0.033160, -0.032352, 0.004581, -0.028335, -0.011976, -0.030335, -0.016279, -0.044635, 0.018961, -0.031429, -0.032280, -0.007870, -0.049753, 0.015269, 0.012114, -0.061564, -0.125598, -0.228144, -0.220672, -0.224792, -0.165259, -0.102422, -0.051713, -0.071218, -0.061103, -0.043678, -0.003041, 0.010492, 0.018285, 0.015490, 0.034521, -0.027878, -0.033017, -0.023685, 0.012960, -0.032718, 0.040195, 0.023083, 0.036129, 0.042083, 0.055360, 0.091629, 0.025951, -0.094581, -0.155765, -0.137664, -0.148806, -0.135908, -0.104630, -0.067548, 0.014486, -0.010555, 0.058674, 0.004691, -0.026710, -0.015717, -0.022107, -0.031037, 0.003459, -0.008668, -0.020270, -0.019192, -0.016304, 0.023208, -0.002732, 0.030924, 0.028715, 0.002224, 0.100582, 0.063131, 0.029619, -0.080669, -0.122975, -0.054604, -0.091045, -0.058839, -0.061809, -0.007083, 0.072895, 0.107448, 0.052351, 0.020531, -0.019265, -0.005755, -0.029845, -0.028269, -0.007895, 0.034025, 0.002734, -0.028132, 0.016048, 0.041645, 0.056271, 0.045029, 0.045922, 0.095747, 0.116869, 0.088558, -0.009624, -0.083637, 0.001317, 0.012563, 0.032163, 0.019118, 0.036547, 0.070636, 0.122451, 0.096961, 0.089529, 0.046947, -0.014567, 0.023073, 0.002786, -0.009053, -0.016032, -0.031921, -0.000211, 0.015267, 0.012621, 0.043878, 0.065576, 0.071440, 0.078941, 0.081830, 0.140047, 0.014283, -0.058289, 0.004634, 0.070282, 0.048794, 0.039489, -0.044224, 0.021804, 0.077992, 0.114436, 0.104772, 0.079841, 0.082958, 0.013606, -0.019797, 0.034314, -0.007458, -0.006609, 0.009049, 0.025399, -0.036346, -0.018494, -0.003381, 0.029129, 0.064467, 0.110009, 0.163125, 0.097525, 0.056385, 0.029925, 0.048092, 0.069325, 0.051241, -0.033377, 0.012762, 0.010677, 0.071069, 0.130239, 0.127819, 0.067387, 0.014873, -0.030793, -0.035985, -0.007967, -0.027728, -0.003614, -0.019281, 0.014256, -0.000360, 0.001177, -0.024838, 0.021747, 0.099543, 0.134905, 0.206654, 0.117568, 0.084773, 0.008041, 0.018384, 0.014698, -0.044791, -0.062701, 0.021726, 0.071221, 0.099121, 0.098210, 0.083595, 0.034673, 0.054171, -0.024207, -0.037528, 0.029577, -0.002880, 0.023983, -0.012494, 0.019823, -0.056523, -0.022963, 0.001722, 0.037571, 0.125998, 0.168678, 0.189375, 0.205090, 0.068327, 0.047218, -0.017084, -0.052724, -0.064517, -0.023371, 0.022193, 0.076439, 0.064360, 0.058109, 0.026645, 0.004013, -0.012536, 0.021195, -0.030167, -0.027634, -0.029077, 0.033400, -0.005240, -0.019683, -0.015656, -0.080460, -0.060229, 0.043782, 0.111933, 0.150350, 0.238674, 0.235592, 0.166950, 0.049359, 0.034524, -0.004025, -0.004034, 0.091965, 0.090778, 0.118356, 0.058748, 0.058934, 0.019304, -0.035409, -0.029631, -0.009918, -0.023149, 0.004407, 0.018859, 0.004151, -0.036020, -0.010859, -0.051985, -0.054908, -0.095856, -0.052847, 0.041273, 0.157245, 0.227734, 0.263464, 0.208512, 0.094968, 0.076053, 0.092179, 0.134295, 0.163561, 0.146090, 0.120279, 0.059710, 0.010855, 0.021044, 0.003238, -0.002716, 0.014538, 0.014302, 0.031166, 0.031068, -0.029135, -0.034617, -0.027832, -0.004898, -0.030841, -0.080685, -0.093992, -0.043031, 0.071375, 0.196141, 0.242013, 0.225516, 0.251485, 0.230242, 0.175110, 0.156454, 0.158066, 0.072009, 0.075458, -0.000328, -0.025957, -0.055131, -0.063628, -0.009346, -0.018965, -0.022015, 0.028468, 0.006622, -0.009584, -0.033598, -0.025854, -0.033978, -0.035834, -0.113617, -0.071570, -0.048524, -0.032247, -0.002684, 0.121963, 0.168035, 0.214698, 0.185337, 0.161237, 0.088294, 0.052652, 0.019893, -0.054672, -0.038364, -0.012896, -0.006943, -0.016887, -0.015920, 0.011555, -0.031774, -0.010757, 0.030977, 0.004596, -0.000773, -0.030837, -0.034222, -0.024399, -0.084734, -0.097026, -0.128389, -0.113866, -0.107880, -0.126710, -0.047233, -0.045896, -0.065796, -0.031848, -0.095078, -0.111063, -0.074006, -0.085105, -0.064117, -0.065280, -0.031546, 0.015807, -0.037440, -0.025563, -0.007931, -0.028265, 0.006685, -0.007097, 0.026937, -0.036446, -0.002739, 0.004340, -0.021030, -0.059359, -0.047367, -0.141429, -0.116242, -0.165657, -0.169305, -0.156584, -0.167848, -0.147320, -0.133699, -0.132967, -0.055000, -0.020537, -0.017365, -0.026048, -0.043294, -0.006643, 0.006737, -0.028558, 0.030307, -0.000940, 0.009754, 0.031507, 0.015498, -0.019469, 0.012213, 0.017559, 0.009186, -0.034638, -0.028352, -0.074345, -0.070868, -0.108209, -0.071516, -0.059743, -0.123889, -0.093805, -0.077655, -0.073960, -0.003590, -0.052952, -0.035195, -0.039581, -0.005491, -0.028998, -0.024836, 0.035413, 0.015951, 0.015152, 0.025328, 0.006171, 0.005795, -0.026846, 0.009787, -0.028914, -0.002920, -0.025044, -0.030452, -0.036191, -0.038629, -0.046213, -0.046660, -0.041197, -0.060218, 0.003599, -0.010148, -0.053943, -0.049585, -0.027451, 0.007771, 0.029105, -0.007350, 0.020303, -0.019568, -0.007419, -0.005541, -0.034771, 0.000186, 0.009452, 0.021768, -0.027642, -0.010856, 0.001133, 0.003082, 0.004570, -0.029113, 0.024138, -0.037518, -0.018907, 0.010678, -0.016395, -0.024294, -0.041493, 0.018564, -0.006376, 0.013049, 0.002689, -0.028656, -0.013723, 0.025142, -0.017550, -0.016467, 0.019583, -0.015479, 0.005830, -0.017362, 0.010993, 0.003633, -0.028348, -0.027089, 0.013112, -0.011753, 0.019478, 0.001720, -0.012397, -0.006489, -0.016591, 0.017048, 0.027560, -0.002080, -0.023796, 0.024876, 0.028238, 0.023768, -0.000997, 0.008584, 0.001697, -0.013685, -0.035372, -0.004365, 0.015447, 0.020833, 0.008494
--  Sum of weights (converted): FFFFFFFFF72FCACE
    );

    constant weights_n7 : weight_array := (
     x"00856A17", x"00B72313", x"80388FA9", x"00BF0C6E", x"80062530", x"80679D79", x"80719CDC", x"80AA82F5", x"80E1568A", x"004305C9", x"010E59DE", x"00299759", x"00278391", x"806E3179", x"8073BF7F", x"805BB759", x"00654515", x"003270F2", x"806B7EE9", x"003953F4", x"80331DF4", x"8013EDC6", x"00CF73C7", x"8079E9F9", x"0110FC70", x"80A006E7", x"010F0EAA", x"006DE977", x"007579D7", x"8042ECE7", x"804FBB47", x"80D6016C", x"81189264", x"00CCD619", x"011B5506", x"0052720F", x"80741B0C", x"003DD88B", x"800D645F", x"8100C016", x"80EF5562", x"0062051D", x"8058738E", x"80489FB8", x"80B3B480", x"007E9722", x"8094C4E2", x"805DFCAB", x"009C223C", x"01192260", x"0104BF3C", x"007322A6", x"000A6496", x"00DBE41E", x"0102ACE8", x"00835903", x"00560112", x"00468C92", x"001DC578", x"00C10AEE", x"00527B35", x"80F6C109", x"80ADD724", x"810D1D38", x"805DFC55", x"0004623E", x"808D399B", x"81238D00", x"80DA76D0", x"005CF6BB", x"8036BE29", x"80520944", x"00105DCE", x"80592ED2", x"80B4AA50", x"8094C69A", x"807F0B49", x"8115DE64", x"81102DE2", x"806F91D4", x"006D8FB5", x"011E197E", x"8007EB32", x"00C7CBEC", x"0060BD82", x"80E90461", x"80925EB9", x"80507ADF", x"80F19368", x"0027A783", x"004130F9", x"80F1BA68", x"805976D0", x"812CAA90", x"00E2A123", x"00571390", x"80D07126", x"0085EB74", x"8137735A", x"006E1F65", x"80F12560", x"8017BC3F", x"0079539D", x"004CF628", x"001F790A", x"803A393C", x"8009999E", x"00F3EECC", x"8061A98B", x"805F0A2B", x"00255836", x"808DF4F7", x"806E9D2E", x"0016DC89", x"00DC08CB", x"005F932A", x"80B65F0C", x"00A5B7E1", x"80811A60", x"00192453", x"804B1BFF", x"00393361", x"811F5980", x"81A080DE", x"81C88C74", x"81E6A0C6", x"82A9DDB4", x"816545CC", x"82A18D50", x"81834E5C", x"82362F14", x"812198BA", x"80F4B6AD", x"80EDEEAB", x"00505FF6", x"81273D84", x"0011465C", x"801F0D5E", x"8099934B", x"00E37B46", x"00B7AA91", x"0058698B", x"0005A04D", x"00A19973", x"808644CD", x"80FB46B7", x"00E73F82", x"80D22633", x"8067756A", x"8107E236", x"80B3E654", x"81555C6C", x"84260500", x"844CF3F0", x"85BA0FC8", x"843BB088", x"83B36D50", x"84C3A4C8", x"8367E7C0", x"831C2DAC", x"8267D6F4", x"8089CC9D", x"81FD7374", x"80B8560D", x"80414508", x"811582BE", x"0072E00D", x"00C2ED26", x"80E86811", x"007131CC", x"800CF2B1", x"0120FFD8", x"8105FB60", x"011FA6F4", x"80305B40", x"01322DB6", x"803854A7", x"004C2552", x"0005178E", x"806302BF", x"81F7AEC6", x"835E556C", x"852FFDF8", x"8641AD38", x"851E7788", x"83B6E590", x"83582844", x"84157190", x"81D06A84", x"813AF23C", x"818A9B10", x"80679161", x"80A3C9F5", x"801F0D1C", x"80D31E2A", x"8025C11C", x"011E6C30", x"00B68270", x"80D794EB", x"0039DF7D", x"0148217A", x"0098C1AB", x"01AD0B4A", x"02F8C674", x"03C5AB68", x"04234CC0", x"02498580", x"01477074", x"01E894F6", x"8059F402", x"8030D9FD", x"8053F29F", x"80C6D783", x"008EBE0C", x"0089B49B", x"8083B72F", x"009D43B8", x"80B7E583", x"813EBB00", x"81FEEB22", x"00102CC8", x"81959D52", x"00C0F91D", x"8067FE0F", x"80361B21", x"003506EA", x"017866C6", x"001B696C", x"0083BCA9", x"02D7ECAC", x"029D88D8", x"03CB9038", x"05561870", x"04702B98", x"05A4EC30", x"042E5F20", x"04DFB5E0", x"048E2C10", x"0410CD78", x"047E48F0", x"065E1758", x"05FC8508", x"045F3ED8", x"03F94C34", x"01742EA2", x"00CC65EE", x"808A416B", x"80DDBE6B", x"80F3474E", x"8077BCA0", x"005BB071", x"00D9CF4D", x"00B6EBE1", x"8061A7A2", x"01889DF4", x"0208B300", x"0260DCB0", x"02CFE898", x"02BD5468", x"035109EC", x"0435BA00", x"036156FC", x"04AA1760", x"03296964", x"0344A0C8", x"04434D10", x"06B40430", x"08589180", x"07B61D50", x"078918B0", x"06AF6660", x"047FC6D8", x"01C70B74", x"01B59014", x"808DBFB3", x"807276AA", x"80481444", x"00A2426E", x"810F8516", x"00DCFD00", x"002E344A", x"011F508A", x"01B0C788", x"0108CAC2", x"01F3C41C", x"026B3ED4", x"03C968F8", x"0265FDFC", x"03298CF4", x"02E60DF0", x"03690978", x"02EC6C00", x"03469F3C", x"0296D5D4", x"03CC0440", x"04F665C0", x"085A7650", x"07F1CFB8", x"06A87B80", x"053C3A98", x"03226998", x"02574360", x"0021DBAC", x"005E28CF", x"81841E00", x"814AE382", x"0055DF9A", x"0112B2FC", x"80684714", x"0135ED16", x"002ED31D", x"005ECB04", x"01C27C44", x"02A4CA14", x"0146CD72", x"02B01418", x"009B49A6", x"00490D27", x"805BEBF9", x"8153063A", x"00B3C1BF", x"8089EAFB", x"80216835", x"01BD1B56", x"05C6C638", x"0638E708", x"05BC1538", x"0395635C", x"03486A6C", x"01C90848", x"016D7186", x"801F7D6F", x"00757164", x"00A6A60A", x"00283B6B", x"8118DCAC", x"003C91AB", x"80C40924", x"00A1A07F", x"00E12584", x"0268A15C", x"0093CA51", x"802D7F34", x"00FC9F30", x"00B70D7A", x"81A62440", x"82C791F8", x"83592194", x"84B76E30", x"85930BB0", x"8414B1D8", x"8089A787", x"024A21A4", x"04B86028", x"03E9BEF0", x"029836E4", x"01D5D054", x"805C1E5B", x"0091AFA6", x"81123520", x"814CAF30", x"802EE03C", x"8076FCEC", x"80B8B301", x"803D99D6", x"8013A50B", x"0098749D", x"00C6C43C", x"00C47968", x"00D9BFAF", x"80D33523", x"003E52A6", x"81299108", x"82E8C904", x"86CD9570", x"86E918C8", x"888DDD80", x"8A7F8610", x"86C39538", x"834373A8", x"017C376E", x"03A51278", x"037E9294", x"03603D48", x"007D2B56", x"01A2EDE8", x"0020677B", x"805FA807", x"81226238", x"809AB1AD", x"011AE6AC", x"00D8B99D", x"00E40963", x"8013EE13", x"80842F98", x"009468BC", x"801956C4", x"8097C947", x"80533C4B", x"80C07005", x"83DD4128", x"863FB670", x"874DA1C8", x"8973AEE0", x"8A9CA3D0", x"8A85B410", x"8797D190", x"829A8BC4", x"028AD24C", x"03BBA610", x"03DFEDDC", x"02BD5494", x"01AAC25A", x"019CFB0A", x"006C27E5", x"812ACB02", x"800DCEC2", x"009EC8D9", x"804CF5E7", x"8036A42F", x"8027A190", x"00B3AC13", x"00FA0FFB", x"80BD1D21", x"00E1EA65", x"0020918E", x"8092A532", x"82CA3750", x"846CCF38", x"84496218", x"868F9350", x"87FF0BD8", x"88901590", x"871A2E88", x"84D3A170", x"00E49B7B", x"0277BC04", x"04613D40", x"044C9D28", x"0259F0CC", x"01DA699E", x"01570514", x"80ACA18C", x"80522E05", x"800B7A4C", x"00E5F738", x"003D8CBC", x"80F91233", x"80555B0C", x"01210A98", x"8026F7FB", x"00E8A9F6", x"0027E2A3", x"002E8030", x"81B3837C", x"8110D342", x"8337F830", x"84BAFBC0", x"8480C238", x"8548A7B0", x"8625F9B8", x"84123F78", x"8012D752", x"028DD7C8", x"02F3C1F8", x"02AC6710", x"01B9BDFC", x"021C9CC8", x"0103F2EE", x"80E02BD4", x"8090ECD1", x"802E6F25", x"814BFBE6", x"00DE6AF5", x"80233F2D", x"80772627", x"002093B7", x"0069A649", x"003CC5D8", x"010A8A2A", x"007DE196", x"80DB36FF", x"817042BA", x"8233257C", x"839EA880", x"84C7BCB8", x"849C5790", x"849EC000", x"8402E070", x"80124CE9", x"0191D478", x"040A7F40", x"02811480", x"01BEF350", x"008A36D3", x"80569191", x"807D9070", x"806A4E7B", x"81312DF6", x"812681B0", x"8015F9F2", x"809CECDC", x"800ED16E", x"0054F6FE", x"00833D16", x"811B06A0", x"006E8E32", x"8087071F", x"8125B920", x"819C256E", x"822D6040", x"82427D04", x"84632E28", x"8397F880", x"83223374", x"83D06250", x"80DCC54F", x"01394AE6", x"03310AA8", x"02835A30", x"805DD5B4", x"809669DD", x"80B98B07", x"824BE350", x"832D5DA0", x"82115140", x"815E676A", x"80BCE32E", x"8096B23D", x"805E04B7", x"80910D0B", x"00BCE597", x"80A54629", x"806132DE", x"00BE1D00", x"80ACF2DA", x"809BB1C0", x"81CBCB38", x"83502AF4", x"82857390", x"84297008", x"84859298", x"83E14E28", x"81E4A484", x"01315754", x"030AED90", x"02550394", x"805AC0CC", x"81330884", x"82543600", x"8237927C", x"83829270", x"842811F0", x"8225CA78", x"82058BAC", x"809E82F1", x"8008546F", x"00505A28", x"009F3718", x"80CD2B52", x"80EE4F1E", x"01122042", x"0101D7FE", x"80A4C18C", x"0080E5E9", x"81182A2C", x"82A2C44C", x"83CF9BE4", x"844F9C50", x"82E36834", x"83A09D54", x"81DF9D14", x"01C3EC0C", x"00DD3F2A", x"01E4E854", x"8025E8F3", x"81923CB2", x"82AE8324", x"83E44558", x"831A1BBC", x"82D036B4", x"82EF0B88", x"827334E4", x"81C0B9FC", x"806A6A00", x"00450024", x"80BB9C17", x"0035E5F1", x"00A8887F", x"00ABEE65", x"80771752", x"0011F343", x"81855392", x"803E9087", x"82CB3724", x"82978C8C", x"835C544C", x"83C1FB60", x"83046EA4", x"816D885A", x"80A47AFD", x"00DA5DBA", x"80BDA919", x"81EA052C", x"81F4B086", x"832C1AC4", x"8377AD4C", x"824DFB78", x"83A24A20", x"82C4E288", x"80D7D40B", x"0031B08C", x"8149D7BE", x"0051C120", x"01206534", x"802F0110", x"80ACA3EE", x"008F85E0", x"009D2B52", x"80416A14", x"813AAAB0", x"80710158", x"81B05D94", x"823B7854", x"80B91F36", x"807E0DFD", x"8059592E", x"8176B8F6", x"0079A1D2", x"00092DA5", x"007D1FAF", x"80A41519", x"8149F84C", x"82C11894", x"819A436A", x"827FF194", x"83131DF8", x"8032DD0B", x"80E92F6C", x"00480955", x"804E3D1F", x"80385710", x"0100FCA6", x"00F2EA66", x"80888CCC", x"00092419", x"00C19F56", x"80012FC8", x"802B8F09", x"01278BC2", x"014525DA", x"0032707F", x"01362606", x"007C1A9B", x"00E1A8FE", x"017E411C", x"001C0892", x"001E4D72", x"00963D15", x"803D0662", x"0134C91A", x"813564D8", x"8214AE48", x"816595E0", x"816C26A4", x"80E14288", x"8071DA27", x"00D4647E", x"8134C95C", x"80BA2D51", x"00359D1E", x"8104753A", x"80E723C8", x"00E02E8C", x"0070356E", x"8053C545", x"008DBB0E", x"00D551E7", x"010725E8", x"02D5B3C8", x"026963CC", x"039269E8", x"023624B4", x"026DBDC4", x"02E70A84", x"039AAF80", x"02A6FD70", x"03B038FC", x"013C2C34", x"00BA5BFB", x"00C3E213", x"8180C2FC", x"81C591CA", x"80CE5907", x"81516056", x"0014B966", x"80493C24", x"805EE4A4", x"00A1C5EA", x"00110599", x"8107C53C", x"81153EBA", x"00B72A7B", x"008827A9", x"00D4BB68", x"80797552", x"00D87B1D", x"02FD1CC0", x"03F01F98", x"0464B3B8", x"050C2D50", x"04136908", x"03A2673C", x"0532C9A0", x"053EC120", x"03CD64A4", x"0311EDE8", x"01F7EC70", x"80386B1C", x"8074FD0C", x"80ABDFF3", x"00383D99", x"807651D1", x"006AB0C2", x"0103BF54", x"803EBC7A", x"8047539F", x"80B7C385", x"80165412", x"810BBDA8", x"00C5C1D7", x"00FC4A3A", x"0052B3DA", x"012D582C", x"00E5EBEB", x"01818AA8", x"025A85D0", x"00F58646", x"0231F31C", x"031CBE24", x"02773628", x"02314894", x"028BFEDC", x"022EFE98", x"01EC15B4", x"00CDCAF2", x"009F4AE2", x"00F5F85C", x"80964D9A", x"007932D4", x"80E6BCEF", x"80B85FA2", x"001E40E5", x"010F5D2C", x"810E31C8", x"007F5970", x"00332B60", x"80EF0FD5", x"80D46D47", x"009367C3", x"8091E6CC", x"00D1353B", x"80C0C571", x"00EC3C98", x"807BF54C", x"00997BB2", x"0089DF86", x"80AC17CE", x"803F9862", x"003DD8E8", x"00A6CB03", x"01250FA8", x"001D897F", x"00B80C24", x"80436EAA", x"8066CC90", x"00C65483", x"804AA2B8", x"80F4C26F", x"000E7D95", x"8029B527", x"00532CA2", x"80953F2E", x"000C99F9"
--  0.016286, 0.022356, -0.006904, 0.023321, -0.000750, -0.012648, -0.013869, -0.020814, -0.027507, 0.008181, 0.033002, 0.005077, 0.004823, -0.013451, -0.014129, -0.011196, 0.012362, 0.006157, -0.013122, 0.006998, -0.006240, -0.002433, 0.025324, -0.014882, 0.033323, -0.019535, 0.033088, 0.013417, 0.014340, -0.008170, -0.009733, -0.026124, -0.034249, 0.025004, 0.034586, 0.010064, -0.014173, 0.007550, -0.001635, -0.031342, -0.029216, 0.011965, -0.010797, -0.008865, -0.021937, 0.015453, -0.018160, -0.011473, 0.019059, 0.034318, 0.031829, 0.014055, 0.001269, 0.026842, 0.031577, 0.016034, 0.010499, 0.008612, 0.003634, 0.023565, 0.010069, -0.030121, -0.021221, -0.032851, -0.011473, 0.000535, -0.017239, -0.035590, -0.026668, 0.011348, -0.006682, -0.010014, 0.001998, -0.010887, -0.022054, -0.018161, -0.015508, -0.033920, -0.033225, -0.013619, 0.013374, 0.034924, -0.000967, 0.024389, 0.011809, -0.028444, -0.017867, -0.009824, -0.029489, 0.004841, 0.007958, -0.029508, -0.010921, -0.036702, 0.027665, 0.010629, -0.025445, 0.016348, -0.038019, 0.013443, -0.029437, -0.002897, 0.014810, 0.009395, 0.003842, -0.007107, -0.001172, 0.029777, -0.011922, -0.011602, 0.004559, -0.017329, -0.013503, 0.002791, 0.026860, 0.011667, -0.022262, 0.020229, -0.015760, 0.003069, -0.009169, 0.006983, -0.035077, -0.050843, -0.055731, -0.059403, -0.083236, -0.043612, -0.082221, -0.047279, -0.069114, -0.035351, -0.029872, -0.029044, 0.009811, -0.036040, 0.002109, -0.003791, -0.018747, 0.027769, 0.022420, 0.010793, 0.000687, 0.019726, -0.016390, -0.030673, 0.028229, -0.025653, -0.012629, -0.032212, -0.021960, -0.041670, -0.129641, -0.134394, -0.178963, -0.132286, -0.115653, -0.148882, -0.106434, -0.097190, -0.075176, -0.016821, -0.062189, -0.022502, -0.007967, -0.033876, 0.014023, 0.023795, -0.028370, 0.013818, -0.001581, 0.035278, -0.031980, 0.035114, -0.005903, 0.037375, -0.006876, 0.009295, 0.000622, -0.012086, -0.061485, -0.105265, -0.162108, -0.195517, -0.159969, -0.116076, -0.104511, -0.127618, -0.056691, -0.038446, -0.048170, -0.012643, -0.019994, -0.003790, -0.025771, -0.004609, 0.034964, 0.022279, -0.026316, 0.007065, 0.040055, 0.018647, 0.052374, 0.092868, 0.117880, 0.129309, 0.071475, 0.039971, 0.059641, -0.010981, -0.005963, -0.010248, -0.024273, 0.017425, 0.016810, -0.016079, 0.019197, -0.022448, -0.038908, -0.062368, 0.001974, -0.049513, 0.023556, -0.012694, -0.006605, 0.006473, 0.045947, 0.003346, 0.016081, 0.088858, 0.081730, 0.118599, 0.166760, 0.138693, 0.176382, 0.130661, 0.152308, 0.142355, 0.127051, 0.140416, 0.198986, 0.187075, 0.136627, 0.124182, 0.045432, 0.024951, -0.016877, -0.027068, -0.029697, -0.014616, 0.011193, 0.026588, 0.022329, -0.011921, 0.047927, 0.063562, 0.074324, 0.087879, 0.085612, 0.103642, 0.131558, 0.105632, 0.145763, 0.098805, 0.102127, 0.133215, 0.209475, 0.260812, 0.240981, 0.235485, 0.208911, 0.140598, 0.055547, 0.053413, -0.017303, -0.013973, -0.008799, 0.019807, -0.033145, 0.026976, 0.005640, 0.035073, 0.052830, 0.032323, 0.061007, 0.075591, 0.118336, 0.074950, 0.098822, 0.090583, 0.106572, 0.091360, 0.102371, 0.080913, 0.118654, 0.155078, 0.261043, 0.248268, 0.208067, 0.163602, 0.097951, 0.073152, 0.004133, 0.011494, -0.047378, -0.040392, 0.010483, 0.033533, -0.012729, 0.037833, 0.005716, 0.011571, 0.054991, 0.082616, 0.039893, 0.083994, 0.018956, 0.008917, -0.011221, -0.041385, 0.021943, -0.016836, -0.004078, 0.054334, 0.180514, 0.194446, 0.179209, 0.111986, 0.102590, 0.055790, 0.044610, -0.003844, 0.014336, 0.020343, 0.004911, -0.034285, 0.007394, -0.023930, 0.019730, 0.027484, 0.075272, 0.018041, -0.005554, 0.030838, 0.022345, -0.051531, -0.086862, -0.104630, -0.147391, -0.174200, -0.127526, -0.016804, 0.071549, 0.147507, 0.122283, 0.081081, 0.057350, -0.011245, 0.017784, -0.033473, -0.040611, -0.005722, -0.014525, -0.022546, -0.007520, -0.002398, 0.018610, 0.024263, 0.023984, 0.026581, -0.025782, 0.007608, -0.036324, -0.090916, -0.212596, -0.215954, -0.267318, -0.328067, -0.211375, -0.101984, 0.046413, 0.113900, 0.109201, 0.105498, 0.015279, 0.051139, 0.003956, -0.011677, -0.035447, -0.018884, 0.034534, 0.026456, 0.027837, -0.002433, -0.016136, 0.018116, -0.003093, -0.018529, -0.010161, -0.023491, -0.120759, -0.195277, -0.228227, -0.295371, -0.331621, -0.328821, -0.237283, -0.081365, 0.079446, 0.116656, 0.121085, 0.085612, 0.052095, 0.050413, 0.013203, -0.036474, -0.001686, 0.019383, -0.009395, -0.006670, -0.004838, 0.021933, 0.030525, -0.023085, 0.027578, 0.003976, -0.017901, -0.087185, -0.138282, -0.133958, -0.205026, -0.249884, -0.267588, -0.221946, -0.150834, 0.027906, 0.077116, 0.136870, 0.134352, 0.073479, 0.057912, 0.041873, -0.021073, -0.010032, -0.001401, 0.028072, 0.007513, -0.030404, -0.010419, 0.035283, -0.004757, 0.028401, 0.004869, 0.005676, -0.053163, -0.033304, -0.100582, -0.147825, -0.140718, -0.165119, -0.192136, -0.127228, -0.002300, 0.079815, 0.092256, 0.083545, 0.053924, 0.065993, 0.031732, -0.027365, -0.017691, -0.005668, -0.040525, 0.027151, -0.004303, -0.014545, 0.003977, 0.012897, 0.007419, 0.032537, 0.015366, -0.026760, -0.044954, -0.068743, -0.113117, -0.149382, -0.144085, -0.144379, -0.125351, -0.002234, 0.049052, 0.126281, 0.078257, 0.054559, 0.016872, -0.010567, -0.015328, -0.012977, -0.037253, -0.035951, -0.002683, -0.019156, -0.001809, 0.010372, 0.016020, -0.034549, 0.013496, -0.016483, -0.035855, -0.050311, -0.068039, -0.070616, -0.137107, -0.112301, -0.097925, -0.119188, -0.026950, 0.038244, 0.099737, 0.078534, -0.011454, -0.018361, -0.022649, -0.071764, -0.099288, -0.064614, -0.042774, -0.023058, -0.018396, -0.011477, -0.017706, 0.023059, -0.020175, -0.011865, 0.023207, -0.021112, -0.019006, -0.056127, -0.103536, -0.078790, -0.130058, -0.141305, -0.121253, -0.059160, 0.037273, 0.095084, 0.072878, -0.011078, -0.037480, -0.072780, -0.069284, -0.109689, -0.129891, -0.067113, -0.063177, -0.019350, -0.001017, 0.009809, 0.019435, -0.025045, -0.029090, 0.033463, 0.031475, -0.020112, 0.015735, -0.034200, -0.082369, -0.119093, -0.134718, -0.090260, -0.113356, -0.058547, 0.055166, 0.027008, 0.059193, -0.004628, -0.049101, -0.083803, -0.121615, -0.096937, -0.087917, -0.091680, -0.076563, -0.054776, -0.012990, 0.008423, -0.022902, 0.006579, 0.020573, 0.020988, -0.014537, 0.002191, -0.047525, -0.007637, -0.087307, -0.081000, -0.105021, -0.117429, -0.094291, -0.044621, -0.020078, 0.026656, -0.023152, -0.059817, -0.061119, -0.099134, -0.108359, -0.072019, -0.113561, -0.086534, -0.026346, 0.006066, -0.040264, 0.009980, 0.035205, -0.005738, -0.021074, 0.017520, 0.019186, -0.007985, -0.038411, -0.013795, -0.052779, -0.069760, -0.022598, -0.015388, -0.010907, -0.045742, 0.014848, 0.001120, 0.015274, -0.020030, -0.040280, -0.086071, -0.050081, -0.078118, -0.096084, -0.006209, -0.028465, 0.008794, -0.009551, -0.006877, 0.031370, 0.029653, -0.016669, 0.001116, 0.023636, -0.000145, -0.005317, 0.036077, 0.039691, 0.006157, 0.037860, 0.015149, 0.027546, 0.046662, 0.003422, 0.003699, 0.018340, -0.007449, 0.037694, -0.037768, -0.065025, -0.043651, -0.044452, -0.027498, -0.013898, 0.025927, -0.037694, -0.022727, 0.006545, -0.031794, -0.028215, 0.027366, 0.013697, -0.010226, 0.017301, 0.026040, 0.032123, 0.088587, 0.075365, 0.111623, 0.069109, 0.075896, 0.090703, 0.112633, 0.082885, 0.115262, 0.038595, 0.022749, 0.023912, -0.046968, -0.055367, -0.025189, -0.041184, 0.002530, -0.008940, -0.011584, 0.019748, 0.002078, -0.032199, -0.033843, 0.022359, 0.016620, 0.025968, -0.014826, 0.026426, 0.093397, 0.123062, 0.137293, 0.157736, 0.127369, 0.113575, 0.162450, 0.163910, 0.118822, 0.095939, 0.061514, -0.006887, -0.014281, -0.020981, 0.006865, -0.014443, 0.013024, 0.031707, -0.007658, -0.008707, -0.022432, -0.002726, -0.032683, 0.024140, 0.030797, 0.010096, 0.036785, 0.028067, 0.047063, 0.073550, 0.029971, 0.068597, 0.097259, 0.077052, 0.068516, 0.079589, 0.068237, 0.060069, 0.025121, 0.019445, 0.030026, -0.018348, 0.014795, -0.028166, -0.022507, 0.003693, 0.033125, -0.032983, 0.015546, 0.006246, -0.029182, -0.025931, 0.017994, -0.017810, 0.025538, -0.023532, 0.028837, -0.015132, 0.018736, 0.016830, -0.021007, -0.007763, 0.007550, 0.020360, 0.035774, 0.003606, 0.022467, -0.008231, -0.012549, 0.024210, -0.009111, -0.029878, 0.001769, -0.005091, 0.010153, -0.018219, 0.001538
--  Sum of weights (converted): FFFFFFFFDD0CEB1A
    );

    constant weights_n8 : weight_array := (
     x"8090565E", x"80B0D1C3", x"0042E139", x"005A6E0E", x"0036203D", x"010E406E", x"001B1F2B", x"0018E11B", x"80263FE4", x"811ADBBA", x"00726E07", x"00E4132E", x"001CEA07", x"80E4C248", x"01063CA6", x"00418639", x"00D39E71", x"007F11B5", x"002E260B", x"80563372", x"003C10C7", x"005E2369", x"8011BCA6", x"80BAE061", x"8099C21A", x"810C27FE", x"80726D72", x"802F2A60", x"00EF493C", x"809C8055", x"811FE1E4", x"00A05C47", x"00FC408E", x"80E4362D", x"80031297", x"005C7FA7", x"00BBB46B", x"803617C0", x"008348F3", x"00DE3F10", x"00A7CB0A", x"008ABAB4", x"00AD9175", x"810A5CC0", x"003936C7", x"00DDCE1F", x"80EA3D72", x"81021C62", x"80F2D37E", x"00590AAE", x"010F285E", x"801A9C4B", x"80744DEC", x"00115080", x"80F13C18", x"0032A582", x"80C059D3", x"80C4EC15", x"80D56BF1", x"8052DE6C", x"00BE5F27", x"003B4F47", x"00CADA91", x"811C91AA", x"80F29FC2", x"00A928BB", x"00D29A3C", x"00DD2195", x"8137BFEC", x"004D3EDC", x"81631FD0", x"809C5561", x"8040A5A7", x"0049BABB", x"808BF4AA", x"81277C7C", x"8133EAE2", x"8083BA03", x"00D6833D", x"007B79AC", x"008F24F2", x"80ED2A37", x"8106E2A4", x"010EB43C", x"00BF1B0A", x"807E1AB5", x"001891D8", x"00D2992C", x"01071280", x"80ED63EB", x"8096B6BE", x"0062B5F7", x"00C36721", x"8003D559", x"806D269D", x"807BC538", x"0055CA8B", x"81C9C0FE", x"809E8864", x"82155158", x"8143808C", x"826E55F0", x"805A9994", x"8185E1EC", x"80788DE4", x"80FEFF6E", x"80002973", x"809332FE", x"80999126", x"807FFEFF", x"00B50CFE", x"0028E300", x"804B5B92", x"00F92E88", x"00397BF4", x"805F1E76", x"801096E7", x"8083E608", x"809E313A", x"80AA7156", x"8035856C", x"81C1C9C6", x"81E19444", x"80630897", x"81626B64", x"80F4B020", x"8017EACF", x"80E1F71C", x"00293E0F", x"8160DD34", x"815EFFEC", x"824F670C", x"80D55557", x"81E249B4", x"800FC3C5", x"80910469", x"808A165D", x"8061E616", x"0072D9B6", x"011F147C", x"004F7C97", x"00B35465", x"80F6DB03", x"804ABA24", x"80BA5359", x"8111490E", x"8056E799", x"8139FED2", x"80E776ED", x"81A87250", x"821ED21C", x"80CFEACC", x"8045377F", x"0205AE44", x"0212EFD4", x"04636348", x"041EC370", x"027B1D34", x"01607F66", x"8074D441", x"008591A7", x"81179916", x"80F68ED6", x"807A57CE", x"00450437", x"8056CD0C", x"008D73F2", x"0095E47A", x"80242640", x"00C1FA0D", x"8101DEFA", x"80B12024", x"8047D3D9", x"8097246A", x"8081B5F6", x"8051E107", x"81BEAAE0", x"0004CAC5", x"002CFDDD", x"019DBD08", x"01F657E8", x"01A3165E", x"0243829C", x"027AD920", x"034E8AF4", x"0373CF14", x"01C95274", x"01E0D1C2", x"00D3C794", x"00966B18", x"001C43C6", x"80AD54BA", x"8030176D", x"00F83E22", x"00F7D60D", x"8063FEA9", x"00F02350", x"00F0441D", x"80FD06DC", x"813A8880", x"80D26F29", x"80AB9FD3", x"8060A06C", x"000CFD97", x"00F3FD0A", x"80013EBC", x"01A97356", x"01017A0C", x"8055EED6", x"80BB1977", x"8060DC82", x"009BD916", x"812FAAC0", x"806CD240", x"80D7EAF2", x"011D6AE6", x"013BFC36", x"0108DF90", x"022B46B4", x"021185FC", x"01863F04", x"001E675B", x"800449BF", x"008BE3D8", x"0062A816", x"80F929B1", x"807984C2", x"00983506", x"80C1DB9E", x"00ABC0B2", x"8020B227", x"02012950", x"00D16381", x"030470F0", x"019938B4", x"0203BC08", x"0186E33C", x"00120A2C", x"82055CB8", x"82598E38", x"831114AC", x"82B72420", x"804BB3B1", x"002B8EFD", x"019508D2", x"02CF8CC0", x"01E720DC", x"024AE7B0", x"01425C78", x"80C8EE92", x"00E96D5C", x"001226A9", x"8113A338", x"8067B445", x"00272714", x"00B5CC89", x"805CCAE0", x"0148BBAC", x"0082EE13", x"0121370A", x"02DF8658", x"0307C980", x"03B3CC40", x"030DC368", x"0045138C", x"817E38C6", x"825F78D4", x"84C56410", x"8303B73C", x"81CEC536", x"81A46FDA", x"01F25C6A", x"01617BD0", x"03D9B7B0", x"02FD50B8", x"02DDEAE4", x"0254EDCC", x"0055ED7D", x"8087205E", x"00860487", x"802F8402", x"01046A0E", x"80E716B5", x"8053C0C5", x"80BD5D4A", x"80060DAA", x"0142594C", x"02211C00", x"031945B8", x"0424A298", x"036AD2A4", x"02327448", x"0217D7DC", x"80C4B25B", x"81B8A51A", x"8338F19C", x"82AB0FC0", x"81FCA6A4", x"801CBAE4", x"01CD08F2", x"028A6F4C", x"0497DA80", x"045ACFC8", x"038ECCB8", x"01028AE4", x"807F96B1", x"00793BFF", x"0107719E", x"802E944E", x"00EA0B6C", x"00C3A4F1", x"004A5A8F", x"802B838F", x"0047CE96", x"01498B64", x"0288682C", x"0351947C", x"02C53AFC", x"0278FB04", x"0287A488", x"0466C050", x"032CC150", x"80A69CE5", x"829D8D58", x"82AE31AC", x"003E9130", x"010EFF4E", x"031C5674", x"02417664", x"04741DB8", x"04004F70", x"0223E6E8", x"00AB5CA3", x"00D35DD9", x"807930F6", x"80773F74", x"006DAD56", x"80E1C172", x"00406AD9", x"801EF8FF", x"00006AF4", x"0048C29B", x"00C9A134", x"003A848B", x"01A3EA98", x"0052F1B4", x"015475BC", x"0178D410", x"0605F0D8", x"0590B5B8", x"02A62614", x"00A8057C", x"005BE1E1", x"8047C618", x"807C65D9", x"0231F36C", x"02D44874", x"020C3538", x"01A1973E", x"00FBACBC", x"00572386", x"00FDB7F6", x"809C02F7", x"81106D1E", x"803060A7", x"80AAF90C", x"80C46EB5", x"80612745", x"80425ADC", x"003A88C7", x"803E1F01", x"804DDDBA", x"80B30EDB", x"818E80A2", x"81AACD9A", x"01DAB1A4", x"053CAB20", x"064564B8", x"02DA711C", x"01F0632A", x"01E49E9C", x"804D00E7", x"805BAB29", x"800DA1F4", x"80A41ACB", x"0075F37E", x"801694B2", x"004D60A8", x"0093BCCD", x"80427C9F", x"00DD33EC", x"000B5017", x"8037C8BA", x"00BEF44A", x"00E0D27E", x"8062AD3B", x"0050B8C2", x"81424314", x"820BC2D4", x"83BF6A98", x"845780D8", x"8448F200", x"83319760", x"018A507E", x"05B82968", x"053654A8", x"04818360", x"033FF450", x"0128AFA2", x"81007A2A", x"83B18804", x"8331F8B8", x"82F0C8BC", x"823FC378", x"817C1066", x"802CC5F5", x"817BAEB4", x"80AB53CA", x"008F62BF", x"00984447", x"804ADC1B", x"80437C6E", x"802BCA72", x"00BE6183", x"006DD17D", x"81D64EBC", x"82304914", x"845D0980", x"84B852D0", x"83E6C3B4", x"824E4190", x"0145A944", x"0646DA38", x"0610A170", x"03814C24", x"012F7592", x"80657FCD", x"823FCC18", x"84931A80", x"84302430", x"833D7BB8", x"81FA8DF4", x"81106DC6", x"819B8A6A", x"8013F4E8", x"000ACEA6", x"001BB0CF", x"80FD4410", x"010EB6DE", x"0081DCAE", x"001AD7AD", x"00522DCF", x"80D10D1E", x"82420D60", x"8284E5C0", x"83574B24", x"80CD2AFB", x"805EC0D2", x"015DD294", x"032E7824", x"05781610", x"04E05F98", x"0075CD83", x"0073E25D", x"800AEC8D", x"83D1FFF0", x"834C45B8", x"84D17940", x"836B5DE8", x"81DD5332", x"80FDD7EF", x"001A6D80", x"006D7944", x"8158C8AE", x"001F8BEF", x"8106AB68", x"00A68C63", x"00560AC2", x"00D82E60", x"000F81F7", x"00133D67", x"818B2392", x"82B27CC4", x"8198E0DE", x"00F3318C", x"01EACD1C", x"05351AC0", x"0555C818", x"053E25D8", x"03888070", x"810756DE", x"8199549E", x"8123D28C", x"81ED4CCA", x"834B95AC", x"820087F4", x"82C859A8", x"81AEFF08", x"827F9664", x"81C54948", x"80009026", x"003DC0BC", x"8091A6F6", x"0065E9D8", x"804CA7FF", x"00A331E0", x"00135640", x"80A024D7", x"80C710F0", x"8274F7F8", x"80899FE7", x"0171FE50", x"03DA372C", x"042BEB90", x"0529C0F8", x"05062380", x"038D49E4", x"8107F5FA", x"8305B2DC", x"8241296C", x"80E6ADFA", x"81D81612", x"82D11CCC", x"81DFA6E4", x"81FF22F4", x"81712AC2", x"80C540F7", x"8155A712", x"8156F070", x"807E6B3A", x"00087546", x"00D682E3", x"006A2AC5", x"80AB0AE3", x"81205998", x"804D68D3", x"8155ECCA", x"8091C225", x"81938580", x"010BB954", x"024604E0", x"03B772B8", x"0315C224", x"01A0A7AE", x"8037CBC7", x"81CD6C1E", x"828C4C1C", x"81BEA3A6", x"81D32270", x"81D32684", x"80014836", x"8169567A", x"81938220", x"814B19B2", x"00878742", x"00CCE07D", x"80EAC992", x"80F99DFC", x"810C9BAC", x"00875B12", x"8075D4A5", x"00DA0435", x"807B18E3", x"006F88E8", x"807FEA02", x"80642BB4", x"00259F78", x"0056542F", x"02077FE4", x"010D8FBE", x"008543DC", x"8046FB9A", x"827F7490", x"8292179C", x"836DBC7C", x"83328B84", x"82EBCC94", x"82BDF34C", x"803D5C9F", x"80121488", x"00DA58A0", x"004D343E", x"0052A709", x"804D0813", x"001DB898", x"8056E161", x"006DF373", x"80852102", x"00B8FD87", x"004FFB6A", x"00877A85", x"806A3DA6", x"80977C91", x"8004442B", x"804938BA", x"015B69BE", x"8058F2AF", x"004FF617", x"80F9B6FE", x"8065399A", x"80422819", x"80314F91", x"81686CB4", x"80A9AC21", x"81ACC218", x"80BC96B8", x"0138B546", x"80917F66", x"00A09E6C", x"80CF202B", x"0095AE49", x"813B6DE6", x"816B37FE", x"806E3949", x"00E6633D", x"0093D090", x"00BC04FF", x"80442D65", x"00F525A9", x"80D49CAA", x"80FCD376", x"822E5910", x"80C102D9", x"80108D09", x"8133671E", x"00DF5863", x"014CF092", x"03EC4A88", x"03E045A4", x"04B253D0", x"0363575C", x"03483404", x"00EE505B", x"0246F058", x"00E9FBE0", x"01F80BDC", x"8058DD2B", x"801EB4E4", x"8070F912", x"80640E4B", x"803245CD", x"00535365", x"01059418", x"00AC5732", x"808D1343", x"0112EA08", x"802FB64B", x"80CA338C", x"803F9A15", x"8178CAD6", x"807A0E56", x"813DF5A4", x"0046476B", x"007AABF6", x"00F2A694", x"044D5578", x"05D33838", x"07291DE8", x"05F346E0", x"0410C518", x"044C2E20", x"03B3045C", x"00FEF647", x"02096CA8", x"80053AAE", x"80B46FF4", x"0072510A", x"800E7B3C", x"80C2ACF9", x"01018930", x"0016EA0E", x"80B78273", x"008636D5", x"0014B52B", x"802F5D12", x"80E3307F", x"80750A2B", x"80333FE7", x"81C9FDEA", x"80D2C07C", x"81EBCF40", x"80B28E52", x"0016676A", x"00824B5A", x"02DB343C", x"0229A700", x"03C9ACE8", x"03256890", x"026AD09C", x"00C385DC", x"00BA2E64", x"011CE8A2", x"01794E1E", x"807E1A12", x"80D0EB22", x"808A2C16", x"80D97908", x"80285E74", x"80D0DE2F", x"00D4225A", x"00CFA9C5", x"80BA293A", x"0101F936", x"00390C94", x"80DC6A44", x"000DE1BF", x"81958B12", x"81815064", x"82254D1C", x"82480E30", x"82003DA0", x"817ECA98", x"81743E2A", x"82664690", x"81E00CD6", x"80A53114", x"007F24E1", x"0001FE18", x"00BA5AC9", x"80B0AFE9", x"0036D832", x"811AD0F4", x"0087D981", x"800E2BB3", x"80190CFB", x"809E5C86", x"80FFE8DD", x"806BB7F5", x"801BA539", x"809B5EEC", x"007A491C", x"803303CE", x"00142F1F", x"81220AFC", x"0033B4B1", x"80BAB5E5", x"811E39B4", x"80CFB216", x"81818A9A", x"8164336C", x"004B15F6", x"006227CE", x"814751D0", x"803150B2", x"80FB089E", x"00C332BE", x"007FE0F1", x"00539983", x"8101B716", x"80994CF1", x"80401B4A", x"8105C824", x"80AB0718", x"004CF7D0", x"80EE2CC8", x"004DD817", x"8006AFA0", x"801817DB", x"80557602", x"809D3C8C", x"81119FFC", x"80C78C42", x"00DBFF5B", x"80171222", x"011AD1D4", x"000C3CCE", x"8028B40C", x"00A986B0", x"811BC99C", x"80BF777D", x"009B081C", x"80573C4F", x"00DCC914", x"8024FE39", x"00C9DF24", x"000B4E8E", x"001CD5C1", x"80F7C8ED", x"8065C853", x"000E96A8", x"0085AD83", x"0038C497", x"803F85A4", x"0001F9AB"
--  -0.017619, -0.021584, 0.008164, 0.011039, 0.006607, 0.032990, 0.003311, 0.003037, -0.004669, -0.034529, 0.013968, 0.027841, 0.003530, -0.027925, 0.032011, 0.007999, 0.025832, 0.015511, 0.005633, -0.010523, 0.007332, 0.011491, -0.002165, -0.022812, -0.018769, -0.032734, -0.013968, -0.005758, 0.029210, -0.019104, -0.035142, 0.019575, 0.030793, -0.027858, -0.000375, 0.011291, 0.022913, -0.006603, 0.016026, 0.027130, 0.020483, 0.016935, 0.021188, -0.032515, 0.006984, 0.027076, -0.028594, -0.031508, -0.029642, 0.010869, 0.033100, -0.003248, -0.014197, 0.002114, -0.029448, 0.006182, -0.023480, -0.024038, -0.026052, -0.010116, 0.023239, 0.007240, 0.024762, -0.034737, -0.029617, 0.020649, 0.025708, 0.026994, -0.038055, 0.009429, -0.043350, -0.019084, -0.007891, 0.009000, -0.017084, -0.036070, -0.037588, -0.016080, 0.026186, 0.015073, 0.017474, -0.028951, -0.032090, 0.033045, 0.023328, -0.015394, 0.002999, 0.025708, 0.032113, -0.028978, -0.018398, 0.012050, 0.023853, -0.000468, -0.013324, -0.015109, 0.010473, -0.055878, -0.019352, -0.065102, -0.039490, -0.075969, -0.011060, -0.047593, -0.014716, -0.031128, -0.000020, -0.017969, -0.018746, -0.015625, 0.022101, 0.004991, -0.009199, 0.030418, 0.007017, -0.011611, -0.002025, -0.016101, -0.019311, -0.020806, -0.006533, -0.054906, -0.058787, -0.012089, -0.043264, -0.029869, -0.002920, -0.027584, 0.005034, -0.043074, -0.042847, -0.072193, -0.026042, -0.058873, -0.001924, -0.017702, -0.016856, -0.011951, 0.014020, 0.035044, 0.009703, 0.021891, -0.030134, -0.009122, -0.022745, -0.033360, -0.010608, -0.038330, -0.028255, -0.051812, -0.066262, -0.025381, -0.008449, 0.063193, 0.064812, 0.137132, 0.128755, 0.077529, 0.043029, -0.014261, 0.016305, -0.034131, -0.030097, -0.014934, 0.008425, -0.010596, 0.017267, 0.018297, -0.004413, 0.023679, -0.031478, -0.021622, -0.008768, -0.018450, -0.015834, -0.009995, -0.054525, 0.000585, 0.005492, 0.050505, 0.061321, 0.051158, 0.070741, 0.077496, 0.103338, 0.107887, 0.055825, 0.058694, 0.025852, 0.018362, 0.003450, -0.021159, -0.005871, 0.030303, 0.030253, -0.012206, 0.029314, 0.029329, -0.030887, -0.038395, -0.025688, -0.020950, -0.011795, 0.001586, 0.029784, -0.000152, 0.051935, 0.031430, -0.010490, -0.022839, -0.011824, 0.019024, -0.037069, -0.013284, -0.026357, 0.034841, 0.038572, 0.032333, 0.067783, 0.064639, 0.047637, 0.003711, -0.000523, 0.017076, 0.012043, -0.030415, -0.014834, 0.018580, -0.023664, 0.020966, -0.003991, 0.062642, 0.025560, 0.094292, 0.049954, 0.062956, 0.047716, 0.002202, -0.063155, -0.073432, -0.095835, -0.084856, -0.009241, 0.005317, 0.049443, 0.087836, 0.059464, 0.071644, 0.039351, -0.024528, 0.028495, 0.002216, -0.033647, -0.012659, 0.004779, 0.022192, -0.011327, 0.040129, 0.015983, 0.035305, 0.089786, 0.094701, 0.115698, 0.095430, 0.008432, -0.046658, -0.074154, -0.149096, -0.094204, -0.056491, -0.051323, 0.060835, 0.043150, 0.120327, 0.093422, 0.089590, 0.072867, 0.010489, -0.016495, 0.016360, -0.005800, 0.031789, -0.028209, -0.010224, -0.023116, -0.000739, 0.039349, 0.066542, 0.096835, 0.129472, 0.106790, 0.068659, 0.065411, -0.024011, -0.053790, -0.100701, -0.083382, -0.062091, -0.003507, 0.056279, 0.079399, 0.143537, 0.136085, 0.111182, 0.031560, -0.015575, 0.014799, 0.032159, -0.005686, 0.028570, 0.023882, 0.009076, -0.005312, 0.008766, 0.040228, 0.079151, 0.103708, 0.086576, 0.077268, 0.079058, 0.137543, 0.099213, -0.020338, -0.081732, -0.083764, 0.007638, 0.033081, 0.097209, 0.070491, 0.139174, 0.125038, 0.066883, 0.020918, 0.025802, -0.014794, -0.014557, 0.013388, -0.027558, 0.007863, -0.003781, 0.000051, 0.008882, 0.024613, 0.007143, 0.051259, 0.010125, 0.041560, 0.046000, 0.188225, 0.173915, 0.082782, 0.020510, 0.011216, -0.008761, -0.015185, 0.068598, 0.088413, 0.063990, 0.050975, 0.030722, 0.010637, 0.030972, -0.019044, -0.033255, -0.005905, -0.020871, -0.023979, -0.011860, -0.008100, 0.007145, -0.007583, -0.009505, -0.021858, -0.048645, -0.052100, 0.057946, 0.163656, 0.195971, 0.089165, 0.060594, 0.059158, -0.009400, -0.011190, -0.001664, -0.020032, 0.014398, -0.002756, 0.009446, 0.018034, -0.008116, 0.027002, 0.001381, -0.006810, 0.023310, 0.027444, -0.012045, 0.009854, -0.039339, -0.063936, -0.117116, -0.135682, -0.133904, -0.099804, 0.048134, 0.178731, 0.162882, 0.140810, 0.101557, 0.036217, -0.031308, -0.115421, -0.099850, -0.091893, -0.070284, -0.046395, -0.005465, -0.046348, -0.020914, 0.017503, 0.018587, -0.009138, -0.008238, -0.005346, 0.023240, 0.013406, -0.057411, -0.068394, -0.136357, -0.147500, -0.121919, -0.072053, 0.039754, 0.196149, 0.189530, 0.109533, 0.037043, -0.012390, -0.070288, -0.142957, -0.130877, -0.101255, -0.061835, -0.033255, -0.050237, -0.002436, 0.001319, 0.003380, -0.030916, 0.033046, 0.015852, 0.003277, 0.010032, -0.025519, -0.070563, -0.078723, -0.104406, -0.025045, -0.011567, 0.042703, 0.099423, 0.170909, 0.152389, 0.014380, 0.014146, -0.001334, -0.119385, -0.103061, -0.150571, -0.106856, -0.058267, -0.030987, 0.003226, 0.013363, -0.042088, 0.003851, -0.032064, 0.020331, 0.010503, 0.026389, 0.001893, 0.002349, -0.048235, -0.084288, -0.049912, 0.029687, 0.059912, 0.162732, 0.166721, 0.163836, 0.110413, -0.032146, -0.049967, -0.035623, -0.060217, -0.102977, -0.062565, -0.086957, -0.052612, -0.078075, -0.055333, -0.000069, 0.007538, -0.017780, 0.012441, -0.009357, 0.019921, 0.002360, -0.019549, -0.024300, -0.076778, -0.016800, 0.045165, 0.120388, 0.130361, 0.161347, 0.156999, 0.110997, -0.032222, -0.094446, -0.070454, -0.028159, -0.057628, -0.088026, -0.058551, -0.062395, -0.045064, -0.024079, -0.041706, -0.041863, -0.015432, 0.001032, 0.026185, 0.012960, -0.020879, -0.035199, -0.009449, -0.041739, -0.017793, -0.049258, 0.032681, 0.071047, 0.116144, 0.096406, 0.050861, -0.006811, -0.056326, -0.079626, -0.054521, -0.057023, -0.057025, -0.000157, -0.044109, -0.049256, -0.040418, 0.016544, 0.025009, -0.028661, -0.030471, -0.032789, 0.016523, -0.014384, 0.026613, -0.015027, 0.013615, -0.015615, -0.012228, 0.004593, 0.010538, 0.063415, 0.032905, 0.016268, -0.008665, -0.078059, -0.080334, -0.107146, -0.099920, -0.091284, -0.085687, -0.007490, -0.002207, 0.026654, 0.009424, 0.010089, -0.009403, 0.003628, -0.010606, 0.013422, -0.016251, 0.022582, 0.009763, 0.016538, -0.012969, -0.018492, -0.000521, -0.008938, 0.042409, -0.010858, 0.009761, -0.030483, -0.012357, -0.008076, -0.006019, -0.043997, -0.020712, -0.052339, -0.023021, 0.038172, -0.017761, 0.019607, -0.025284, 0.018272, -0.038505, -0.044338, -0.013455, 0.028123, 0.018044, 0.022952, -0.008322, 0.029925, -0.025954, -0.030863, -0.068158, -0.023561, -0.002020, -0.037525, 0.027264, 0.040642, 0.122594, 0.121127, 0.146768, 0.105877, 0.102564, 0.029091, 0.071160, 0.028562, 0.061529, -0.010848, -0.003748, -0.013791, -0.012214, -0.006137, 0.010172, 0.031931, 0.021038, -0.017221, 0.033559, -0.005824, -0.024683, -0.007764, -0.045995, -0.014899, -0.038813, 0.008579, 0.014975, 0.029620, 0.134440, 0.182034, 0.223769, 0.185947, 0.127047, 0.134299, 0.115603, 0.031123, 0.063650, -0.000638, -0.022026, 0.013955, -0.001768, -0.023764, 0.031437, 0.002797, -0.022401, 0.016384, 0.002528, -0.005782, -0.027733, -0.014287, -0.006256, -0.055907, -0.025727, -0.060035, -0.021796, 0.002735, 0.015905, 0.089258, 0.067585, 0.118369, 0.098316, 0.075539, 0.023868, 0.022727, 0.034779, 0.046058, -0.015393, -0.025503, -0.016867, -0.026547, -0.004928, -0.025497, 0.025895, 0.025350, -0.022725, 0.031491, 0.006964, -0.026906, 0.001695, -0.049505, -0.047035, -0.067053, -0.071296, -0.062529, -0.046727, -0.045440, -0.074985, -0.058600, -0.020165, 0.015521, 0.000243, 0.022748, -0.021568, 0.006695, -0.034523, 0.016583, -0.001730, -0.003058, -0.019331, -0.031239, -0.013149, -0.003375, -0.018966, 0.014927, -0.006227, 0.002464, -0.035406, 0.006312, -0.022792, -0.034940, -0.025353, -0.047063, -0.043482, 0.009166, 0.011982, -0.039956, -0.006020, -0.030644, 0.023828, 0.015610, 0.010205, -0.031459, -0.018713, -0.007826, -0.031956, -0.020877, 0.009396, -0.029074, 0.009502, -0.000816, -0.002941, -0.010432, -0.019194, -0.033401, -0.024359, 0.026855, -0.002816, 0.034524, 0.001494, -0.004969, 0.020694, -0.034642, -0.023372, 0.018925, -0.010649, 0.026951, -0.004516, 0.024643, 0.001380, 0.003520, -0.030247, -0.012425, 0.001781, 0.016318, 0.006930, -0.007754, 0.000241
--  Sum of weights (converted): 000000005DB9074C
    );

    constant weights_n9 : weight_array := (
     x"00FB80AC", x"00C329EA", x"0063D4B0", x"80D2D96E", x"80625FD9", x"00BACA25", x"01075DAA", x"808A5037", x"007C50A5", x"80448217", x"00B998A7", x"802BF620", x"80E8B8E1", x"81226564", x"800B77FD", x"00563B01", x"80AC781E", x"00E62FFE", x"008AC67C", x"00B06DFA", x"0086CBA5", x"811A2E9E", x"8035A4D9", x"0097F8F7", x"0090D47E", x"810A3396", x"80A5D705", x"00D54037", x"80F23AC8", x"00DDBD43", x"8038727E", x"001576C9", x"008EAEEE", x"004EB930", x"80BC19E1", x"005DCDE0", x"80FD34BC", x"80967227", x"8036D9F2", x"80405117", x"00CD02EB", x"80A692A2", x"00EF2240", x"008149F4", x"0056661A", x"00CA543A", x"80CB3F97", x"80FE5163", x"00094BC6", x"008F82F5", x"00933C40", x"000C0A59", x"0117D134", x"0067F232", x"007E6B00", x"808DCE4C", x"00593ED5", x"806D8402", x"80EC5A0C", x"80BE6B16", x"80B1037F", x"802C3D8C", x"807B7FC4", x"0108BD4E", x"00729D09", x"80FE588E", x"80099BCB", x"00DC82C7", x"8039D95D", x"800C49BA", x"000B5CB2", x"80A55580", x"810065AC", x"80A8A501", x"807DD9AF", x"00C02B08", x"8102AF46", x"001BB2DF", x"80764B4B", x"8020FF16", x"801A8CBD", x"8071B73B", x"004382A7", x"0045253E", x"80A802E7", x"00B3C2F7", x"0107EA54", x"80797F37", x"003B4FB1", x"806DA70A", x"00C442DB", x"8022D9B0", x"811B5F14", x"001CEE91", x"00AEC439", x"8060928C", x"80CEC8D1", x"80B6138D", x"802ECE22", x"000DC5D7", x"812F56DA", x"802DE721", x"0004F0A2", x"008927FD", x"00806862", x"81200E16", x"810682D2", x"80FBC87D", x"00B4D15A", x"80950761", x"00A18085", x"802B9009", x"80788E25", x"00DC27D4", x"80388437", x"809E3146", x"802E7F1C", x"80C25292", x"812EC4CC", x"805F8BF3", x"8064A3E0", x"813A21AC", x"00238F18", x"8179F6FA", x"82077DD8", x"81546C2C", x"828736C4", x"832DBD7C", x"82BDBFA8", x"83B4DF8C", x"810C4BEA", x"815C36E6", x"80CB8B70", x"81AC6042", x"006407BB", x"812AE08A", x"807C183C", x"80C1DE55", x"8095E813", x"003E59D4", x"81222598", x"811E6BB0", x"0042CA3A", x"005E8883", x"80066656", x"80997CDA", x"80B96100", x"80E823D8", x"816ECE6E", x"828B12E4", x"8173833C", x"825968B8", x"84082D00", x"843C9A40", x"85AB6360", x"864BE788", x"85B2B340", x"860E9C98", x"85075478", x"848E22B0", x"83A5DA54", x"82597870", x"829468B8", x"82419E08", x"0044F388", x"8021F642", x"00AA90D4", x"00DC0733", x"007FF71E", x"806407C4", x"8037668D", x"8018F85B", x"801C1CF2", x"807E0A29", x"81F67926", x"827BA2C4", x"81DF57F6", x"8315F684", x"8395B31C", x"819B8ADC", x"81A61110", x"80031126", x"030C3B98", x"020A5FA8", x"01984E16", x"016793F0", x"81077212", x"82D360BC", x"82213054", x"831F785C", x"8402A6E8", x"82F99778", x"8178EAEE", x"80806211", x"80F62148", x"8070FF39", x"0062E345", x"81126BEE", x"811944A8", x"0026E6AD", x"80488B21", x"8242F278", x"831193D4", x"821B5C48", x"82668060", x"83D89AD8", x"811EFDF4", x"0093D935", x"03B56970", x"05ACD9A8", x"093101A0", x"0B4E79E0", x"096F1AB0", x"0489A4E0", x"0293A0D0", x"008B81D5", x"82B87ADC", x"83F064B4", x"845ACA00", x"83677C60", x"8222A294", x"8159CC66", x"812C144E", x"00B40C61", x"011DA07E", x"00EEDC15", x"009C4FEE", x"0028FAA2", x"814313F8", x"82734950", x"82DE5DB4", x"828D66DC", x"827FD5FC", x"81FD064E", x"810049CC", x"011168D0", x"031DF098", x"0540DE78", x"061531F0", x"06434F98", x"043C96C8", x"0263E208", x"000A585C", x"8042192A", x"82723114", x"81E10D24", x"83E90C40", x"833325CC", x"8088E807", x"80F00ED6", x"805E35FC", x"0093CA49", x"80FD4962", x"804CFA8E", x"80335532", x"804E7E2C", x"8121C87A", x"8207E060", x"8242AFBC", x"814ED0BE", x"003CDC6E", x"00210620", x"02431430", x"03A7F938", x"018204D4", x"02323964", x"0168C46A", x"808D5DF0", x"003C58EE", x"006F5DF6", x"00DBF5B1", x"008F6E7F", x"804890E7", x"80B84B0A", x"82AF6FDC", x"81D0C186", x"8037BED6", x"80FC61E0", x"0022FD3C", x"80994E49", x"006AB319", x"0053486F", x"00ABE60C", x"806B26B3", x"801FD725", x"006E6FF5", x"00A6C548", x"00029A3E", x"030391E8", x"023680E0", x"044A9D48", x"024DDD44", x"00D4FBD2", x"823A2ED0", x"83AF552C", x"81D68DF4", x"817A99E2", x"0002070C", x"015542B0", x"02A63064", x"021F57D8", x"00AA6F5B", x"80409BF9", x"807C4E60", x"805F02CC", x"00929CA8", x"0093C33A", x"809A8905", x"802D718F", x"007CF62E", x"00B83B1B", x"8140A7F4", x"80A2501C", x"00920C6F", x"03477C48", x"0457BA80", x"038155A0", x"03C8923C", x"03CF3498", x"016DCED2", x"821C13E8", x"83BDEB48", x"82A83800", x"80845826", x"015DE1EC", x"03AB7B38", x"03D746BC", x"05D78838", x"035B785C", x"01AFFC7C", x"016246B2", x"80798A9C", x"8163F362", x"006E36CF", x"8080F6EA", x"0119F3B8", x"8055759E", x"80E3034F", x"80F9CDCA", x"80147E58", x"0086986D", x"02FC9FB4", x"033ABACC", x"032B9EA4", x"04422038", x"032EA240", x"028EF0A8", x"802D6F26", x"83251480", x"81C96D52", x"00588BC4", x"023188CC", x"03B692CC", x"06657658", x"0609C2B8", x"06C7C638", x"0397A998", x"030AEF20", x"8034B8D7", x"81304D1C", x"005F2FCD", x"00C39067", x"806F48F4", x"00FFEB90", x"0020F07F", x"0066594E", x"802464A1", x"80385DFD", x"00BFFB9D", x"0177E578", x"03E45C28", x"0410A6D0", x"04ABE708", x"01EA5F98", x"02183EE0", x"802FFE03", x"8076E7C8", x"0059FC50", x"0371AE84", x"04889AF0", x"067889B0", x"0621F5D0", x"07068390", x"05850E68", x"01998AB8", x"01DD9BC4", x"004D1503", x"81C418AC", x"81A1FDAC", x"8023E6E7", x"00E037A9", x"00540F59", x"0028AC20", x"80144E97", x"812B9AA4", x"00E03E67", x"01D01614", x"00FB8EAA", x"01F7D67E", x"037ECA98", x"023D9498", x"01595F48", x"015770C2", x"0057ACA4", x"0118E2C6", x"0035784A", x"0184C240", x"02C8A120", x"06572A48", x"073AAD60", x"04B4A940", x"019AF1C2", x"8045E51E", x"81D3F310", x"8119726E", x"8077531E", x"816E2B56", x"80FB0AC0", x"00D43940", x"002743CE", x"808A15E5", x"00BD5D93", x"80F54515", x"806F6D2F", x"005CE462", x"00DCDB52", x"011AF462", x"01D7C514", x"019B0F14", x"02088958", x"0139B1D2", x"00583957", x"008D6FD2", x"805A3262", x"80D69C7F", x"001D7F54", x"05766438", x"04A238B8", x"017F1974", x"81282806", x"812DE172", x"81BFEB16", x"83516A3C", x"817E5E70", x"804AEB80", x"0009FC42", x"80122765", x"808AF180", x"80CE86DF", x"8120A0AC", x"800BD194", x"806AD0E4", x"008C960A", x"80721646", x"009862C7", x"80A03806", x"026732F4", x"018FDACA", x"029CF6FC", x"015946EA", x"00638D32", x"8193C4AE", x"817C4ACA", x"006058A8", x"04AC4458", x"037FD100", x"8157AB1C", x"8210206C", x"82DFE13C", x"82A4DDF4", x"81845AC0", x"81CE3C7A", x"816C416C", x"80CE7744", x"0017C488", x"802BC0F9", x"80D18AD3", x"0007DD16", x"009EA2B4", x"800CC4E5", x"00781CE7", x"813BBE0A", x"804781F6", x"80A0262E", x"80958ECD", x"0103C418", x"016F96B4", x"803143CB", x"814D85C4", x"81D600E6", x"8219AE48", x"02687610", x"02839964", x"00190583", x"8191C1DA", x"8228F768", x"82027624", x"821D5558", x"83291A80", x"826EF8BC", x"806510B6", x"00DD051F", x"00EF3CDE", x"00726410", x"0115FC28", x"80867051", x"8012D2A8", x"8122876A", x"8144F6F0", x"8218ABD8", x"82DF7E8C", x"81DF73DC", x"81F0BB28", x"81AB852C", x"812F1508", x"831370E0", x"832D2FF8", x"8180934E", x"80FDF505", x"01CD5212", x"009E503B", x"81D4A144", x"81BFF9EA", x"81DCF31E", x"81D82E52", x"82B35910", x"8184274C", x"80910E79", x"0009F49F", x"8050FAC6", x"81112EAA", x"011E21D6", x"00516B73", x"010216DC", x"0059CEAE", x"803D916A", x"80190341", x"80D0F8AE", x"8264CC6C", x"82FB4388", x"84074C40", x"83F4C0C8", x"8468B978", x"84FCC2E0", x"832535C0", x"81656CEC", x"003562AA", x"80987475", x"8142B68E", x"82E0A278", x"8161BB1A", x"824032A4", x"826D93B0", x"817B67AA", x"828A3618", x"809F6F54", x"80FAC714", x"802289BB", x"8074812E", x"00EC854F", x"80D9762E", x"00348111", x"80087EAE", x"815EE19E", x"00319F8D", x"811D896A", x"835122E4", x"84C8FF30", x"84587D60", x"84F6C070", x"868D3F40", x"862DDA90", x"85788EA0", x"81A9B8BC", x"82256250", x"82AC9A80", x"8212CFE0", x"81CB8992", x"81BEF366", x"80D27978", x"800F5BB0", x"812F7B3E", x"80BAA878", x"809CCFFB", x"80DB8382", x"002F7CEB", x"809B5F16", x"00A94D8D", x"80C9CF89", x"80EF863E", x"8042B934", x"009E1556", x"8167A162", x"8180962C", x"8241D808", x"83F09A88", x"840AC2A8", x"845587C0", x"84F465F0", x"8561BB58", x"84BF8588", x"839C6BB0", x"82EC8FB0", x"83A4A364", x"840313D8", x"829A6EA8", x"8263E774", x"80967F4B", x"81123A06", x"8088A4B8", x"80A65B3E", x"0091948C", x"8101393A", x"80773926", x"003B13BD", x"80526D52", x"80050256", x"00C5B837", x"001FFE23", x"8000E964", x"800AFA16", x"818079BE", x"82320670", x"824209A0", x"8349C980", x"83239E2C", x"840D4E78", x"82781C70", x"823547F8", x"831D3CE4", x"83D3D1C0", x"83937D4C", x"83EF96F4", x"82B5FF14", x"80F22EC0", x"803D0DD1", x"00E101C7", x"800C059E", x"014958D8", x"805DE82A", x"80789955", x"00C52C8B", x"8039482A", x"0053B282", x"8033F957", x"80CEEA73", x"800FF5C5", x"00744C5F", x"0085CEE2", x"0059ECA2", x"810D4DF4", x"80C0252E", x"81569442", x"81E98AC4", x"81C461DA", x"81F50C9C", x"81AFC4A8", x"82911358", x"8232DB8C", x"83329F88", x"825389F4", x"8048AC66", x"80414251", x"01E04B12", x"025A7A8C", x"01795BD8", x"00B4C118", x"00746000", x"00B26E44", x"80DF1F68", x"804ED96D", x"80B240B3", x"8108A164", x"80D155EC", x"80BCA715", x"00D5701F", x"009DFF61", x"80D6439E", x"80FCE911", x"011371B0", x"008410D3", x"00FD25F1", x"010F388E", x"005C7626", x"80124E1B", x"006ABD2C", x"8198B8FA", x"80CD9EB7", x"019EF0EE", x"020B8034", x"02F48880", x"03603EA4", x"01E71B16", x"012B0738", x"005F8B07", x"806C711A", x"0004C2FB", x"00F5F865", x"80137E5B", x"00A07455", x"80918057", x"001D0750", x"80DB5343", x"80174DB2", x"003F37AA", x"804D0D21", x"01641360", x"01096EAA", x"01CFF04E", x"0305C5DC", x"0333495C", x"02D8B2FC", x"03A00EC8", x"040A2BB8", x"01BA50A6", x"029A5514", x"0404A1D0", x"038E6D34", x"02B2BE10", x"02694E60", x"01D606CE", x"01F98120", x"016998D2", x"002A3FC6", x"80E120CE", x"002961B8", x"005019A5", x"806E5C22", x"0064E22B", x"8077837C", x"00627E17", x"00D21C13", x"00A1D555", x"8001D1F4", x"0144A1FA", x"00116A2D", x"80C3DDF0", x"013EABB4", x"019FBE24", x"013B8216", x"01E3B61E", x"018E87C0", x"0190C5FC", x"01669C78", x"000438A0", x"00FDBCF6", x"008A7D10", x"014EF06C", x"8027EE15", x"0076E309", x"0089FE5D", x"80670149", x"80756614", x"80BDDC93", x"00508D80", x"80F595B1", x"803C0D74", x"001045F9", x"00537955", x"80FB2BEA", x"003AF092", x"8073DFE3", x"80236849", x"80D48978", x"80E82862", x"00227973", x"002B5B3C", x"00EE01BF", x"00FF8F71", x"00B16AC9", x"00552575", x"009E781E", x"0056EA7A", x"8133A520", x"00C7AF0C", x"00286A18", x"803C05DB", x"805163D1", x"00EBD2C7", x"00CBFCF5", x"801B2D54", x"806D5E39", x"809D4C5E", x"00A8A9E7"
--  0.030701, 0.023824, 0.012186, -0.025738, -0.012009, 0.022801, 0.032149, -0.016884, 0.015175, -0.008363, 0.022656, -0.005366, -0.028408, -0.035449, -0.001400, 0.010526, -0.021053, 0.028099, 0.016940, 0.021537, 0.016455, -0.034446, -0.006548, 0.018551, 0.017679, -0.032495, -0.020244, 0.026032, -0.029569, 0.027068, -0.006891, 0.002620, 0.017417, 0.009610, -0.022962, 0.011451, -0.030909, -0.018365, -0.006696, -0.007851, 0.025026, -0.020334, 0.029191, 0.015782, 0.010547, 0.024698, -0.024811, -0.031045, 0.001135, 0.017518, 0.017973, 0.001470, 0.034157, 0.012689, 0.015432, -0.017310, 0.010894, -0.013369, -0.028852, -0.023244, -0.021608, -0.005400, -0.015076, 0.032317, 0.013991, -0.031048, -0.001173, 0.026918, -0.007062, -0.001500, 0.001387, -0.020182, -0.031298, -0.020586, -0.015363, 0.023458, -0.031578, 0.003381, -0.014440, -0.004028, -0.003241, -0.013881, 0.008241, 0.008441, -0.020509, 0.021944, 0.032216, -0.014831, 0.007240, -0.013385, 0.023958, -0.004254, -0.034591, 0.003532, 0.021334, -0.011789, -0.025242, -0.022226, -0.005714, 0.001681, -0.037029, -0.005603, 0.000603, 0.016743, 0.015675, -0.035163, -0.032045, -0.030735, 0.022072, -0.018192, 0.019715, -0.005318, -0.014716, 0.026874, -0.006899, -0.019311, -0.005676, -0.023721, -0.036959, -0.011663, -0.012285, -0.038346, 0.004341, -0.046138, -0.063414, -0.041555, -0.079006, -0.099334, -0.085663, -0.115829, -0.032751, -0.042507, -0.024847, -0.052292, 0.012211, -0.036484, -0.015148, -0.023666, -0.018299, 0.007611, -0.035418, -0.034963, 0.008153, 0.011540, -0.000781, -0.018736, -0.022629, -0.028337, -0.044776, -0.079477, -0.045351, -0.073414, -0.125998, -0.132398, -0.177171, -0.196766, -0.178064, -0.189284, -0.157145, -0.142351, -0.113996, -0.073422, -0.080616, -0.070510, 0.008417, -0.004146, 0.020821, 0.026859, 0.015621, -0.012211, -0.006763, -0.003048, -0.003432, -0.015386, -0.061337, -0.077592, -0.058514, -0.096431, -0.112024, -0.050237, -0.051522, -0.000374, 0.095243, 0.063766, 0.049842, 0.043894, -0.032159, -0.088303, -0.066551, -0.097592, -0.125324, -0.092968, -0.046010, -0.015672, -0.030045, -0.013794, 0.012071, -0.033499, -0.034334, 0.004749, -0.008855, -0.070672, -0.095896, -0.065840, -0.075012, -0.120191, -0.035033, 0.018048, 0.115895, 0.177350, 0.287232, 0.353330, 0.294813, 0.141802, 0.080521, 0.017030, -0.085020, -0.123095, -0.136083, -0.106383, -0.066728, -0.042212, -0.036631, 0.021979, 0.034867, 0.029158, 0.019081, 0.005002, -0.039438, -0.076573, -0.089644, -0.079761, -0.078105, -0.062137, -0.031285, 0.033375, 0.097405, 0.164169, 0.190087, 0.195717, 0.132396, 0.074693, 0.001263, -0.008069, -0.076439, -0.058722, -0.122198, -0.099994, -0.016712, -0.029304, -0.011500, 0.018041, -0.030919, -0.009397, -0.006266, -0.009582, -0.035374, -0.063461, -0.070640, -0.040871, 0.007429, 0.004031, 0.070688, 0.114255, 0.047121, 0.068631, 0.044039, -0.017257, 0.007367, 0.013595, 0.026851, 0.017509, -0.008858, -0.022497, -0.083916, -0.056733, -0.006805, -0.030808, 0.004271, -0.018714, 0.013025, 0.010166, 0.020984, -0.013080, -0.003887, 0.013481, 0.020358, 0.000318, 0.094186, 0.069153, 0.134108, 0.072005, 0.025999, -0.069602, -0.115153, -0.057441, -0.046216, 0.000248, 0.041658, 0.082787, 0.066326, 0.020805, -0.007887, -0.015174, -0.011598, 0.017897, 0.018037, -0.018864, -0.005547, 0.015254, 0.022489, -0.039143, -0.019814, 0.017828, 0.102476, 0.135709, 0.109538, 0.118234, 0.119044, 0.044654, -0.065927, -0.116933, -0.083035, -0.016155, 0.042710, 0.114683, 0.120029, 0.182560, 0.104916, 0.052733, 0.043247, -0.014837, -0.043451, 0.013454, -0.015743, 0.034418, -0.010432, -0.027712, -0.030494, -0.002502, 0.016430, 0.093338, 0.100919, 0.099075, 0.133072, 0.099443, 0.079949, -0.005546, -0.098276, -0.055838, 0.010809, 0.068547, 0.116037, 0.199886, 0.188691, 0.211887, 0.112263, 0.095085, -0.006436, -0.037146, 0.011619, 0.023873, -0.013585, 0.031240, 0.004021, 0.012494, -0.004443, -0.006881, 0.023435, 0.045886, 0.121626, 0.127033, 0.145984, 0.059860, 0.065460, -0.005858, -0.014515, 0.010985, 0.107627, 0.141675, 0.202214, 0.191646, 0.219545, 0.172492, 0.049993, 0.058302, 0.009409, -0.055188, -0.051024, -0.004383, 0.027370, 0.010261, 0.004965, -0.002479, -0.036573, 0.027374, 0.056651, 0.030708, 0.061504, 0.109227, 0.070017, 0.042160, 0.041924, 0.010702, 0.034288, 0.006527, 0.047456, 0.086991, 0.198140, 0.225913, 0.147053, 0.050164, -0.008532, -0.057123, -0.034356, -0.014566, -0.044698, -0.030645, 0.025906, 0.004793, -0.016856, 0.023116, -0.029940, -0.013602, 0.011339, 0.026960, 0.034540, 0.057589, 0.050178, 0.063542, 0.038293, 0.010770, 0.017265, -0.011010, -0.026198, 0.003601, 0.170702, 0.144802, 0.046765, -0.036152, -0.036851, -0.054678, -0.103688, -0.046676, -0.009145, 0.001219, -0.002216, -0.016961, -0.025211, -0.035233, -0.001443, -0.013039, 0.017161, -0.013927, 0.018602, -0.019558, 0.075098, 0.048810, 0.081661, 0.042148, 0.012152, -0.049288, -0.046422, 0.011761, 0.146029, 0.109353, -0.041952, -0.064469, -0.089829, -0.082625, -0.047407, -0.056425, -0.044465, -0.025203, 0.002901, -0.005341, -0.025579, 0.000960, 0.019365, -0.001559, 0.014662, -0.038543, -0.008729, -0.019549, -0.018257, 0.031710, 0.044872, -0.006014, -0.040713, -0.057373, -0.065635, 0.075252, 0.078564, 0.003054, -0.049043, -0.067501, -0.062800, -0.066081, -0.098768, -0.076046, -0.012337, 0.026980, 0.029204, 0.013964, 0.033934, -0.016411, -0.002298, -0.035465, -0.039669, -0.065512, -0.089782, -0.058527, -0.060636, -0.052188, -0.036997, -0.096123, -0.099266, -0.046945, -0.031001, 0.056314, 0.019325, -0.057206, -0.054685, -0.058221, -0.057639, -0.084393, -0.047382, -0.017707, 0.001215, -0.009885, -0.033347, 0.034928, 0.009939, 0.031505, 0.010963, -0.007516, -0.003053, -0.025509, -0.074805, -0.093172, -0.125891, -0.123627, -0.137784, -0.155855, -0.098292, -0.043631, 0.006517, -0.018610, -0.039394, -0.089921, -0.043180, -0.070337, -0.075876, -0.046314, -0.079371, -0.019462, -0.030613, -0.004216, -0.014222, 0.028872, -0.026546, 0.006409, -0.001037, -0.042832, 0.006058, -0.034856, -0.103654, -0.149536, -0.135802, -0.155121, -0.204742, -0.193097, -0.170966, -0.051968, -0.067063, -0.083570, -0.064796, -0.056096, -0.054559, -0.025693, -0.001875, -0.037046, -0.022785, -0.019142, -0.026796, 0.005797, -0.018966, 0.020667, -0.024635, -0.029239, -0.008145, 0.019297, -0.043900, -0.046947, -0.070538, -0.123121, -0.126314, -0.135441, -0.154834, -0.168180, -0.148379, -0.112844, -0.091377, -0.113847, -0.125376, -0.081352, -0.074695, -0.018371, -0.033475, -0.016680, -0.020307, 0.017771, -0.031399, -0.014554, 0.007212, -0.010062, -0.000611, 0.024136, 0.003905, -0.000111, -0.001340, -0.046933, -0.068607, -0.070561, -0.102757, -0.098098, -0.126624, -0.077162, -0.069004, -0.097319, -0.119607, -0.111754, -0.122997, -0.084716, -0.029563, -0.007453, 0.027467, -0.001468, 0.040203, -0.011463, -0.014722, 0.024069, -0.006992, 0.010217, -0.006344, -0.025258, -0.001948, 0.014197, 0.016334, 0.010977, -0.032874, -0.023455, -0.041819, -0.059759, -0.055222, -0.061163, -0.052706, -0.080209, -0.068708, -0.099930, -0.072698, -0.008871, -0.007966, 0.058630, 0.073545, 0.046064, 0.022065, 0.014206, 0.021781, -0.027237, -0.009625, -0.021759, -0.032304, -0.025554, -0.023029, 0.026054, 0.019287, -0.026155, -0.030873, 0.033624, 0.016121, 0.030902, 0.033108, 0.011287, -0.002235, 0.013030, -0.049893, -0.025100, 0.050652, 0.063904, 0.092350, 0.105499, 0.059461, 0.036502, 0.011663, -0.013238, 0.000581, 0.030026, -0.002380, 0.019587, -0.017761, 0.003544, -0.026773, -0.002845, 0.007717, -0.009406, 0.043466, 0.032401, 0.056633, 0.094455, 0.100011, 0.088953, 0.113288, 0.126242, 0.053994, 0.081339, 0.125565, 0.111136, 0.084319, 0.075355, 0.057376, 0.061707, 0.044140, 0.005157, -0.027481, 0.005051, 0.009778, -0.013472, 0.012315, -0.014589, 0.012023, 0.025648, 0.019755, -0.000222, 0.039628, 0.002126, -0.023910, 0.038900, 0.050750, 0.038514, 0.059047, 0.048649, 0.048923, 0.043776, 0.000515, 0.030974, 0.016905, 0.040886, -0.004874, 0.014513, 0.016845, -0.012574, -0.014331, -0.023176, 0.009833, -0.029979, -0.007331, 0.001986, 0.010190, -0.030661, 0.007195, -0.014145, -0.004322, -0.025944, -0.028340, 0.004208, 0.005293, 0.029054, 0.031196, 0.021657, 0.010394, 0.019344, 0.010610, -0.037554, 0.024375, 0.004933, -0.007327, -0.009935, 0.028787, 0.024901, -0.003318, -0.013351, -0.019201, 0.020589
--  Sum of weights (converted): FFFFFFFF918181A6
    );

    attribute rom_style : string;
    attribute rom_style of weights_n0 : constant is "block";
    attribute rom_style of weights_n1 : constant is "block";
    attribute rom_style of weights_n2 : constant is "block";
    attribute rom_style of weights_n3 : constant is "block";
    attribute rom_style of weights_n4 : constant is "block";
    attribute rom_style of weights_n5 : constant is "block";
    attribute rom_style of weights_n6 : constant is "block";
    attribute rom_style of weights_n7 : constant is "block";
    attribute rom_style of weights_n8 : constant is "block";
    attribute rom_style of weights_n9 : constant is "block";

begin

    read_n0 : process(clk) is
    begin
        if rising_edge(clk) then
            dout((1*DATA_WIDTH-1) downto (0*DATA_WIDTH)) <= weights_n0(to_integer(unsigned(addr)));
        end if;
    end process read_n0;

    read_n1 : process(clk) is
    begin
        if rising_edge(clk) then
            dout((2*DATA_WIDTH-1) downto (1*DATA_WIDTH)) <= weights_n1(to_integer(unsigned(addr)));
        end if;
    end process read_n1;

    read_n2 : process(clk) is
    begin
        if rising_edge(clk) then
            dout((3*DATA_WIDTH-1) downto (2*DATA_WIDTH)) <= weights_n2(to_integer(unsigned(addr)));
        end if;
    end process read_n2;

    read_n3 : process(clk) is
    begin
        if rising_edge(clk) then
            dout((4*DATA_WIDTH-1) downto (3*DATA_WIDTH)) <= weights_n3(to_integer(unsigned(addr)));
        end if;
    end process read_n3;

    read_n4 : process(clk) is
    begin
        if rising_edge(clk) then
            dout((5*DATA_WIDTH-1) downto (4*DATA_WIDTH)) <= weights_n4(to_integer(unsigned(addr)));
        end if;
    end process read_n4;

    read_n5 : process(clk) is
    begin
        if rising_edge(clk) then
            dout((6*DATA_WIDTH-1) downto (5*DATA_WIDTH)) <= weights_n5(to_integer(unsigned(addr)));
        end if;
    end process read_n5;

    read_n6 : process(clk) is
    begin
        if rising_edge(clk) then
            dout((7*DATA_WIDTH-1) downto (6*DATA_WIDTH)) <= weights_n6(to_integer(unsigned(addr)));
        end if;
    end process read_n6;

    read_n7 : process(clk) is
    begin
        if rising_edge(clk) then
            dout((8*DATA_WIDTH-1) downto (7*DATA_WIDTH)) <= weights_n7(to_integer(unsigned(addr)));
        end if;
    end process read_n7;

    read_n8 : process(clk) is
    begin
        if rising_edge(clk) then
            dout((9*DATA_WIDTH-1) downto (8*DATA_WIDTH)) <= weights_n8(to_integer(unsigned(addr)));
        end if;
    end process read_n8;

    read_n9 : process(clk) is
    begin
        if rising_edge(clk) then
            dout((10*DATA_WIDTH-1) downto (9*DATA_WIDTH)) <= weights_n9(to_integer(unsigned(addr)));
        end if;
    end process read_n9;

end rtl;